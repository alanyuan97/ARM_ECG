module rom_input(EN,data_add,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I74x);
	input EN;
	input [9:0]data_add;
	output reg [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I74x;
	always@(EN)
		begin
		case(data_add)
			10'b0000000000:begin
				I0x <= 8175;
				I1x <= 4726;
				I2x <= 2908;
				I3x <= 1327;
				I4x <= 1310;
				I5x <= 1433;
				I6x <= 1449;
				I7x <= 1384;
				I8x <= 1425;
				I9x <= 1384;
				I10x <= 1368;
				I11x <= 1400;
				I12x <= 1400;
				I13x <= 1449;
				I14x <= 1425;
				I15x <= 1433;
				I16x <= 1507;
				I17x <= 1540;
				I18x <= 1638;
				I19x <= 1662;
				I20x <= 1712;
				I21x <= 1835;
				I22x <= 1916;
				I23x <= 2072;
				I24x <= 2154;
				I25x <= 2260;
				I26x <= 2424;
				I27x <= 2498;
				I28x <= 2629;
				I29x <= 2654;
				I30x <= 2703;
				I31x <= 2760;
				I32x <= 2670;
				I33x <= 2564;
				I34x <= 2285;
				I35x <= 2072;
				I36x <= 1908;
				I37x <= 1712;
				I38x <= 1638;
				I39x <= 1507;
				I40x <= 1441;
				I41x <= 1441;
				I42x <= 1409;
				I43x <= 1441;
				I44x <= 1392;
				I45x <= 1376;
				I46x <= 1400;
				I47x <= 1384;
				I48x <= 1449;
				I49x <= 1409;
				I50x <= 1400;
				I51x <= 1409;
				I52x <= 1400;
				I53x <= 1458;
				I54x <= 1409;
				I55x <= 1400;
				I56x <= 1425;
				I57x <= 1400;
				I58x <= 1449;
				I59x <= 1392;
				I60x <= 1359;
				I61x <= 1359;
				I62x <= 1343;
				I63x <= 1376;
				I64x <= 1318;
				I65x <= 1302;
				I66x <= 1327;
				I67x <= 1310;
				I68x <= 1359;
				I69x <= 1318;
				I70x <= 1335;
				I71x <= 1482;
				I72x <= 1548;
				I73x <= 1654;
				I74x <= 1581;
			end

			10'b0000000001:begin
				I0x <= 8192;
				I1x <= 3407;
				I2x <= 1957;
				I3x <= 478;
				I4x <= 667;
				I5x <= 1441;
				I6x <= 1916;
				I7x <= 1957;
				I8x <= 2048;
				I9x <= 1982;
				I10x <= 2015;
				I11x <= 2064;
				I12x <= 2023;
				I13x <= 2170;
				I14x <= 2228;
				I15x <= 2260;
				I16x <= 2277;
				I17x <= 2269;
				I18x <= 2416;
				I19x <= 2449;
				I20x <= 2441;
				I21x <= 2523;
				I22x <= 2670;
				I23x <= 2752;
				I24x <= 2801;
				I25x <= 2908;
				I26x <= 2949;
				I27x <= 3080;
				I28x <= 3104;
				I29x <= 3112;
				I30x <= 3260;
				I31x <= 3358;
				I32x <= 3399;
				I33x <= 3342;
				I34x <= 3162;
				I35x <= 2998;
				I36x <= 2490;
				I37x <= 2342;
				I38x <= 2228;
				I39x <= 1933;
				I40x <= 1785;
				I41x <= 1818;
				I42x <= 1843;
				I43x <= 1875;
				I44x <= 1843;
				I45x <= 1802;
				I46x <= 1916;
				I47x <= 1892;
				I48x <= 1859;
				I49x <= 1851;
				I50x <= 1933;
				I51x <= 1916;
				I52x <= 1875;
				I53x <= 1957;
				I54x <= 1925;
				I55x <= 1875;
				I56x <= 1818;
				I57x <= 1687;
				I58x <= 1695;
				I59x <= 1802;
				I60x <= 1679;
				I61x <= 1720;
				I62x <= 1728;
				I63x <= 1679;
				I64x <= 1818;
				I65x <= 1736;
				I66x <= 1695;
				I67x <= 1662;
				I68x <= 1703;
				I69x <= 1695;
				I70x <= 1900;
				I71x <= 2236;
				I72x <= 2498;
				I73x <= 2662;
				I74x <= 2883;
			end

			10'b0000000010:begin
				I0x <= 8192;
				I1x <= 6881;
				I2x <= 3522;
				I3x <= 1441;
				I4x <= 0;
				I5x <= 412;
				I6x <= 966;
				I7x <= 901;
				I8x <= 909;
				I9x <= 909;
				I10x <= 909;
				I11x <= 958;
				I12x <= 950;
				I13x <= 958;
				I14x <= 1040;
				I15x <= 1146;
				I16x <= 1155;
				I17x <= 1122;
				I18x <= 1228;
				I19x <= 1302;
				I20x <= 1277;
				I21x <= 1384;
				I22x <= 1466;
				I23x <= 1540;
				I24x <= 1589;
				I25x <= 1654;
				I26x <= 1875;
				I27x <= 2056;
				I28x <= 2220;
				I29x <= 2465;
				I30x <= 2613;
				I31x <= 2826;
				I32x <= 2957;
				I33x <= 3055;
				I34x <= 3121;
				I35x <= 3088;
				I36x <= 2981;
				I37x <= 2768;
				I38x <= 2498;
				I39x <= 2211;
				I40x <= 1949;
				I41x <= 1630;
				I42x <= 1474;
				I43x <= 1376;
				I44x <= 1261;
				I45x <= 1146;
				I46x <= 1073;
				I47x <= 1056;
				I48x <= 1048;
				I49x <= 925;
				I50x <= 950;
				I51x <= 991;
				I52x <= 991;
				I53x <= 991;
				I54x <= 933;
				I55x <= 909;
				I56x <= 999;
				I57x <= 1007;
				I58x <= 1015;
				I59x <= 1007;
				I60x <= 1032;
				I61x <= 1024;
				I62x <= 1015;
				I63x <= 1024;
				I64x <= 1056;
				I65x <= 991;
				I66x <= 1015;
				I67x <= 1032;
				I68x <= 917;
				I69x <= 966;
				I70x <= 983;
				I71x <= 991;
				I72x <= 917;
				I73x <= 942;
				I74x <= 933;
			end

			10'b0000000011:begin
				I0x <= 7667;
				I1x <= 6447;
				I2x <= 3588;
				I3x <= 1622;
				I4x <= 50;
				I5x <= 0;
				I6x <= 424;
				I7x <= 694;
				I8x <= 670;
				I9x <= 697;
				I10x <= 717;
				I11x <= 738;
				I12x <= 774;
				I13x <= 792;
				I14x <= 810;
				I15x <= 843;
				I16x <= 942;
				I17x <= 991;
				I18x <= 1040;
				I19x <= 1056;
				I20x <= 1163;
				I21x <= 1245;
				I22x <= 1286;
				I23x <= 1351;
				I24x <= 1449;
				I25x <= 1548;
				I26x <= 1703;
				I27x <= 1867;
				I28x <= 2048;
				I29x <= 2220;
				I30x <= 2433;
				I31x <= 2637;
				I32x <= 2826;
				I33x <= 2957;
				I34x <= 3006;
				I35x <= 3014;
				I36x <= 2949;
				I37x <= 2744;
				I38x <= 2514;
				I39x <= 2228;
				I40x <= 1925;
				I41x <= 1703;
				I42x <= 1531;
				I43x <= 1368;
				I44x <= 1253;
				I45x <= 1155;
				I46x <= 1089;
				I47x <= 1056;
				I48x <= 1015;
				I49x <= 1015;
				I50x <= 999;
				I51x <= 958;
				I52x <= 958;
				I53x <= 950;
				I54x <= 991;
				I55x <= 1024;
				I56x <= 1024;
				I57x <= 1015;
				I58x <= 1048;
				I59x <= 1040;
				I60x <= 1073;
				I61x <= 1064;
				I62x <= 1040;
				I63x <= 1024;
				I64x <= 1040;
				I65x <= 1081;
				I66x <= 1056;
				I67x <= 1056;
				I68x <= 1040;
				I69x <= 999;
				I70x <= 991;
				I71x <= 966;
				I72x <= 974;
				I73x <= 983;
				I74x <= 966;
			end

			10'b0000000100:begin
				I0x <= 7708;
				I1x <= 4603;
				I2x <= 2940;
				I3x <= 1802;
				I4x <= 1925;
				I5x <= 2023;
				I6x <= 2007;
				I7x <= 1957;
				I8x <= 1982;
				I9x <= 1990;
				I10x <= 2007;
				I11x <= 2023;
				I12x <= 2048;
				I13x <= 2088;
				I14x <= 2097;
				I15x <= 2146;
				I16x <= 2162;
				I17x <= 2211;
				I18x <= 2293;
				I19x <= 2334;
				I20x <= 2400;
				I21x <= 2473;
				I22x <= 2547;
				I23x <= 2686;
				I24x <= 2809;
				I25x <= 2924;
				I26x <= 3039;
				I27x <= 3145;
				I28x <= 3227;
				I29x <= 3268;
				I30x <= 3309;
				I31x <= 3301;
				I32x <= 3227;
				I33x <= 3022;
				I34x <= 2777;
				I35x <= 2547;
				I36x <= 2351;
				I37x <= 2187;
				I38x <= 2080;
				I39x <= 2031;
				I40x <= 1949;
				I41x <= 1933;
				I42x <= 1933;
				I43x <= 1941;
				I44x <= 1933;
				I45x <= 1908;
				I46x <= 1900;
				I47x <= 1900;
				I48x <= 1925;
				I49x <= 1925;
				I50x <= 1908;
				I51x <= 1900;
				I52x <= 1892;
				I53x <= 1875;
				I54x <= 1908;
				I55x <= 1900;
				I56x <= 1875;
				I57x <= 1892;
				I58x <= 1875;
				I59x <= 1875;
				I60x <= 1859;
				I61x <= 1884;
				I62x <= 1859;
				I63x <= 1859;
				I64x <= 1843;
				I65x <= 1859;
				I66x <= 1843;
				I67x <= 1818;
				I68x <= 1818;
				I69x <= 1810;
				I70x <= 1794;
				I71x <= 1777;
				I72x <= 1785;
				I73x <= 1777;
				I74x <= 1777;
			end

			10'b0000000101:begin
				I0x <= 8192;
				I1x <= 7192;
				I2x <= 4161;
				I3x <= 1728;
				I4x <= 1277;
				I5x <= 1236;
				I6x <= 1310;
				I7x <= 1433;
				I8x <= 1400;
				I9x <= 1400;
				I10x <= 1531;
				I11x <= 1302;
				I12x <= 1359;
				I13x <= 1523;
				I14x <= 1376;
				I15x <= 1392;
				I16x <= 1466;
				I17x <= 1597;
				I18x <= 1818;
				I19x <= 1622;
				I20x <= 1925;
				I21x <= 1851;
				I22x <= 2211;
				I23x <= 2285;
				I24x <= 2359;
				I25x <= 2662;
				I26x <= 2875;
				I27x <= 3055;
				I28x <= 3301;
				I29x <= 3571;
				I30x <= 4005;
				I31x <= 3964;
				I32x <= 4038;
				I33x <= 4317;
				I34x <= 4218;
				I35x <= 4366;
				I36x <= 3907;
				I37x <= 3416;
				I38x <= 3047;
				I39x <= 2719;
				I40x <= 2383;
				I41x <= 2539;
				I42x <= 2023;
				I43x <= 1916;
				I44x <= 1818;
				I45x <= 1785;
				I46x <= 1638;
				I47x <= 1540;
				I48x <= 1753;
				I49x <= 1622;
				I50x <= 1638;
				I51x <= 1679;
				I52x <= 1622;
				I53x <= 1605;
				I54x <= 1622;
				I55x <= 1654;
				I56x <= 1802;
				I57x <= 1777;
				I58x <= 1703;
				I59x <= 1671;
				I60x <= 1613;
				I61x <= 1687;
				I62x <= 2105;
				I63x <= 1605;
				I64x <= 1564;
				I65x <= 1589;
				I66x <= 1540;
				I67x <= 1564;
				I68x <= 1794;
				I69x <= 1736;
				I70x <= 1392;
				I71x <= 1622;
				I72x <= 1376;
				I73x <= 1433;
				I74x <= 1835;
			end

			10'b0000000110:begin
				I0x <= 8126;
				I1x <= 7741;
				I2x <= 1753;
				I3x <= 257;
				I4x <= 0;
				I5x <= 295;
				I6x <= 1032;
				I7x <= 1204;
				I8x <= 1212;
				I9x <= 1236;
				I10x <= 1228;
				I11x <= 1236;
				I12x <= 1269;
				I13x <= 1335;
				I14x <= 1327;
				I15x <= 1335;
				I16x <= 1359;
				I17x <= 1441;
				I18x <= 1474;
				I19x <= 1449;
				I20x <= 1474;
				I21x <= 1556;
				I22x <= 1662;
				I23x <= 1744;
				I24x <= 1802;
				I25x <= 1941;
				I26x <= 2023;
				I27x <= 2080;
				I28x <= 2195;
				I29x <= 2441;
				I30x <= 2670;
				I31x <= 2899;
				I32x <= 3186;
				I33x <= 3424;
				I34x <= 3653;
				I35x <= 3784;
				I36x <= 3932;
				I37x <= 4038;
				I38x <= 3956;
				I39x <= 3751;
				I40x <= 3342;
				I41x <= 2908;
				I42x <= 2441;
				I43x <= 2056;
				I44x <= 1695;
				I45x <= 1376;
				I46x <= 1212;
				I47x <= 991;
				I48x <= 950;
				I49x <= 876;
				I50x <= 876;
				I51x <= 876;
				I52x <= 819;
				I53x <= 876;
				I54x <= 909;
				I55x <= 999;
				I56x <= 1024;
				I57x <= 1040;
				I58x <= 1015;
				I59x <= 1015;
				I60x <= 1015;
				I61x <= 1040;
				I62x <= 1081;
				I63x <= 1064;
				I64x <= 1081;
				I65x <= 1024;
				I66x <= 999;
				I67x <= 983;
				I68x <= 942;
				I69x <= 884;
				I70x <= 884;
				I71x <= 843;
				I72x <= 819;
				I73x <= 795;
				I74x <= 753;
			end

			10'b0000000111:begin
				I0x <= 7954;
				I1x <= 6291;
				I2x <= 1703;
				I3x <= 0;
				I4x <= 217;
				I5x <= 1269;
				I6x <= 1802;
				I7x <= 1982;
				I8x <= 2072;
				I9x <= 2129;
				I10x <= 2154;
				I11x <= 2228;
				I12x <= 2269;
				I13x <= 2318;
				I14x <= 2318;
				I15x <= 2326;
				I16x <= 2342;
				I17x <= 2408;
				I18x <= 2457;
				I19x <= 2547;
				I20x <= 2564;
				I21x <= 2719;
				I22x <= 2867;
				I23x <= 2990;
				I24x <= 3121;
				I25x <= 3252;
				I26x <= 3416;
				I27x <= 3620;
				I28x <= 3883;
				I29x <= 4128;
				I30x <= 4382;
				I31x <= 4595;
				I32x <= 4775;
				I33x <= 4833;
				I34x <= 4734;
				I35x <= 4489;
				I36x <= 4112;
				I37x <= 3751;
				I38x <= 3399;
				I39x <= 3039;
				I40x <= 2744;
				I41x <= 2588;
				I42x <= 2473;
				I43x <= 2359;
				I44x <= 2375;
				I45x <= 2334;
				I46x <= 2293;
				I47x <= 2285;
				I48x <= 2203;
				I49x <= 2146;
				I50x <= 2113;
				I51x <= 2097;
				I52x <= 2113;
				I53x <= 2080;
				I54x <= 2097;
				I55x <= 2080;
				I56x <= 2138;
				I57x <= 2105;
				I58x <= 2121;
				I59x <= 2138;
				I60x <= 2146;
				I61x <= 2097;
				I62x <= 2080;
				I63x <= 2064;
				I64x <= 2064;
				I65x <= 2039;
				I66x <= 2048;
				I67x <= 2056;
				I68x <= 2072;
				I69x <= 2072;
				I70x <= 2105;
				I71x <= 2072;
				I72x <= 2048;
				I73x <= 2056;
				I74x <= 2121;
			end

			10'b0000001000:begin
				I0x <= 8019;
				I1x <= 7626;
				I2x <= 3956;
				I3x <= 0;
				I4x <= 1105;
				I5x <= 2260;
				I6x <= 3637;
				I7x <= 3063;
				I8x <= 2473;
				I9x <= 2744;
				I10x <= 2793;
				I11x <= 2662;
				I12x <= 2990;
				I13x <= 2859;
				I14x <= 3014;
				I15x <= 3178;
				I16x <= 3203;
				I17x <= 3383;
				I18x <= 3375;
				I19x <= 3497;
				I20x <= 3776;
				I21x <= 3833;
				I22x <= 4358;
				I23x <= 4407;
				I24x <= 5087;
				I25x <= 5054;
				I26x <= 5152;
				I27x <= 5603;
				I28x <= 5701;
				I29x <= 5668;
				I30x <= 5660;
				I31x <= 5611;
				I32x <= 5611;
				I33x <= 5177;
				I34x <= 4947;
				I35x <= 4300;
				I36x <= 4161;
				I37x <= 3866;
				I38x <= 3440;
				I39x <= 3629;
				I40x <= 3252;
				I41x <= 3129;
				I42x <= 3186;
				I43x <= 3121;
				I44x <= 3309;
				I45x <= 3145;
				I46x <= 3104;
				I47x <= 3252;
				I48x <= 3153;
				I49x <= 3276;
				I50x <= 3153;
				I51x <= 3219;
				I52x <= 3252;
				I53x <= 3219;
				I54x <= 3252;
				I55x <= 3211;
				I56x <= 3104;
				I57x <= 3801;
				I58x <= 3981;
				I59x <= 4210;
				I60x <= 4407;
				I61x <= 4620;
				I62x <= 4726;
				I63x <= 4751;
				I64x <= 4718;
				I65x <= 5062;
				I66x <= 4448;
				I67x <= 4186;
				I68x <= 3538;
				I69x <= 3211;
				I70x <= 2891;
				I71x <= 2727;
				I72x <= 2760;
				I73x <= 2572;
				I74x <= 2629;
			end

			10'b0000001001:begin
				I0x <= 7774;
				I1x <= 7184;
				I2x <= 3948;
				I3x <= 1712;
				I4x <= 364;
				I5x <= 1736;
				I6x <= 2670;
				I7x <= 2809;
				I8x <= 2924;
				I9x <= 3014;
				I10x <= 3129;
				I11x <= 3211;
				I12x <= 3252;
				I13x <= 3268;
				I14x <= 3260;
				I15x <= 3203;
				I16x <= 3301;
				I17x <= 3432;
				I18x <= 3481;
				I19x <= 3538;
				I20x <= 3825;
				I21x <= 3760;
				I22x <= 3956;
				I23x <= 4235;
				I24x <= 4521;
				I25x <= 4808;
				I26x <= 5136;
				I27x <= 5505;
				I28x <= 5816;
				I29x <= 6094;
				I30x <= 6250;
				I31x <= 6381;
				I32x <= 6250;
				I33x <= 5881;
				I34x <= 5365;
				I35x <= 4767;
				I36x <= 4177;
				I37x <= 3653;
				I38x <= 3268;
				I39x <= 2891;
				I40x <= 2826;
				I41x <= 2736;
				I42x <= 2662;
				I43x <= 2588;
				I44x <= 2555;
				I45x <= 2605;
				I46x <= 2588;
				I47x <= 2498;
				I48x <= 2490;
				I49x <= 2531;
				I50x <= 2514;
				I51x <= 2547;
				I52x <= 2506;
				I53x <= 2572;
				I54x <= 2605;
				I55x <= 2621;
				I56x <= 2646;
				I57x <= 2629;
				I58x <= 2703;
				I59x <= 2678;
				I60x <= 2686;
				I61x <= 2686;
				I62x <= 2621;
				I63x <= 2588;
				I64x <= 2596;
				I65x <= 2588;
				I66x <= 2555;
				I67x <= 2588;
				I68x <= 2498;
				I69x <= 2564;
				I70x <= 2416;
				I71x <= 2449;
				I72x <= 2301;
				I73x <= 2342;
				I74x <= 2318;
			end

		endcase
	end
endmodule
