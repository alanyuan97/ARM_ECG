module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [7:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [7:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 8'b10101001;
	I1x = 8'b11010001;
	I2x = 8'b10001011;
	I3x = 8'b11110001;
	I4x = 8'b11010011;
	I5x = 8'b01110111;
	I6x = 8'b00101010;
	I7x = 8'b10101111;
	I8x = 8'b01111011;
	I9x = 8'b01100001;
	I10x = 8'b11111010;
	I11x = 8'b10000010;
	I12x = 8'b00111101;
	I13x = 8'b00010111;
	I14x = 8'b10111001;
	I15x = 8'b00010001;
	I16x = 8'b01000001;
	I17x = 8'b01100100;
	I18x = 8'b00010110;
	I19x = 8'b10101100;
	I20x = 8'b11010101;
	I21x = 8'b01111010;
	I22x = 8'b10001111;
	I23x = 8'b00011011;
	I24x = 8'b11001010;
	I25x = 8'b01000000;
	I26x = 8'b01001100;
	I27x = 8'b01010111;
	I28x = 8'b11100100;
	I29x = 8'b01111100;
	I30x = 8'b10010000;
	I31x = 8'b00110111;
	I32x = 8'b10110111;
	I33x = 8'b01101110;
	I34x = 8'b10111010;
	I35x = 8'b11000001;
	I36x = 8'b00110111;
	I37x = 8'b00111010;
	I38x = 8'b01010011;
	I39x = 8'b01011110;
	I40x = 8'b10111001;
	I41x = 8'b10111000;
	I42x = 8'b00000111;
	I43x = 8'b11111100;
	I44x = 8'b10011000;
	I45x = 8'b10111111;
	I46x = 8'b00110001;
	I47x = 8'b01000110;
	I48x = 8'b01010001;
	I49x = 8'b10110101;
	I50x = 8'b10110100;
	I51x = 8'b00011111;
	I52x = 8'b01001001;
	I53x = 8'b00111110;
	I54x = 8'b11101010;
	I55x = 8'b00111111;
	I56x = 8'b00100011;
	I57x = 8'b11000100;
	I58x = 8'b00010101;
	I59x = 8'b00011001;
	I60x = 8'b01110100;
	I61x = 8'b01001100;
	I62x = 8'b11111001;
	I63x = 8'b11011111;
	I64x = 8'b00111110;
	I65x = 8'b00111100;
	I66x = 8'b10001100;
	I67x = 8'b11000100;
	I68x = 8'b11101011;
	I69x = 8'b11111001;
	I70x = 8'b10111011;
	I71x = 8'b10110001;
	I72x = 8'b01001011;
	I73x = 8'b00000011;
	I74x = 8'b10100010;
	I75x = 8'b10100011;
	I76x = 8'b10000000;
	I77x = 8'b10101011;
	I78x = 8'b10111100;
	I79x = 8'b11001001;
	I80x = 8'b10000110;
	I81x = 8'b00101101;
	I82x = 8'b01100010;
	I83x = 8'b00110001;
	I84x = 8'b01110001;
	I85x = 8'b00000010;
	I86x = 8'b01110001;
	I87x = 8'b00010100;
	I88x = 8'b01100111;
	I89x = 8'b00011010;
	I90x = 8'b11001000;
	I91x = 8'b11101011;
	I92x = 8'b00111100;
	I93x = 8'b01111111;
	I94x = 8'b11000100;
	I95x = 8'b11111100;
	I96x = 8'b11011101;
	I97x = 8'b11110101;
	I98x = 8'b11011000;
	I99x = 8'b00111001;
	I100x = 8'b10110110;
	I101x = 8'b11100011;
	I102x = 8'b11011001;
	I103x = 8'b10011010;
	I104x = 8'b10001001;
	I105x = 8'b01100010;
	I106x = 8'b11111101;
	I107x = 8'b01010101;
	I108x = 8'b01100111;
	I109x = 8'b00000011;
	I110x = 8'b11001110;
	I111x = 8'b11001010;
	I112x = 8'b10111110;
	I113x = 8'b10111110;
	I114x = 8'b11001010;
	I115x = 8'b10001010;
	I116x = 8'b11011010;
	I117x = 8'b10001000;
	I118x = 8'b10011011;
	I119x = 8'b00110001;
	I120x = 8'b10110101;
	I121x = 8'b01011101;
	I122x = 8'b00000010;
	I123x = 8'b11111101;
	I124x = 8'b01000100;
	I125x = 8'b00111111;
	I126x = 8'b00110010;
	I127x = 8'b01001011;
	I128x = 8'b10000001;
	I129x = 8'b10010101;
	I130x = 8'b01010011;
	I131x = 8'b10000111;
	I132x = 8'b11011011;
	I133x = 8'b00001101;
	I134x = 8'b01011000;
	I135x = 8'b10100000;
	I136x = 8'b11101101;
	I137x = 8'b01110101;
	I138x = 8'b00111100;
	I139x = 8'b11010011;
	I140x = 8'b01010100;
	I141x = 8'b00000110;
	I142x = 8'b00011101;
	I143x = 8'b10111011;
	I144x = 8'b11000010;
	I145x = 8'b00111010;
	I146x = 8'b01100110;
	I147x = 8'b10111100;
	I148x = 8'b11110000;
	I149x = 8'b00100010;
	I150x = 8'b00111000;
	I151x = 8'b00011111;
	I152x = 8'b10101110;
	I153x = 8'b01101100;
	I154x = 8'b01110001;
	I155x = 8'b11011010;
	I156x = 8'b01100011;
	I157x = 8'b00001110;
	I158x = 8'b01111010;
	I159x = 8'b10011100;
	I160x = 8'b11011100;
	I161x = 8'b11011100;
	I162x = 8'b01111101;
	I163x = 8'b00100011;
	I164x = 8'b10111001;
	I165x = 8'b01100100;
	I166x = 8'b00101001;
	I167x = 8'b00011011;
	I168x = 8'b00110011;
	I169x = 8'b10101101;
	I170x = 8'b11001010;
	I171x = 8'b11101101;
	I172x = 8'b01010100;
	I173x = 8'b01111001;
	I174x = 8'b11000011;
	I175x = 8'b10110010;
	I176x = 8'b10000111;
	I177x = 8'b00000100;
	I178x = 8'b00001000;
	I179x = 8'b01010100;
	I180x = 8'b10111111;
	I181x = 8'b00101000;
	I182x = 8'b11000000;
	I183x = 8'b01010111;
	I184x = 8'b10110011;
	I185x = 8'b11001000;
	I186x = 8'b01110100;
	end
endmodule
[0.26100502 1.89132649 0.73922447 0.         0.        ] ['00100001', '01111111', '01011110', '00000000', '00000000']
