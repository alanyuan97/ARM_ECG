module node_1_1(clk,reset,N1x,A0x,A1x,A2x,A3x,A4x,A5x,A6x,A7x,A8x,A9x,A10x,A11x,A12x,A13x,A14x,A15x,A16x,A17x,A18x,A19x,A20x,A21x,A22x,A23x,A24x,A25x,A26x,A27x,A28x,A29x,A30x,A31x,A32x,A33x,A34x,A35x,A36x,A37x,A38x,A39x,A40x,A41x,A42x,A43x,A44x,A45x,A46x,A47x,A48x,A49x,A50x,A51x,A52x,A53x,A54x,A55x,A56x,A57x,A58x,A59x,A60x,A61x,A62x,A63x,A64x,A65x,A66x,A67x,A68x,A69x,A70x,A71x,A72x,A73x,A74x,A75x,A76x,A77x,A78x,A79x,A80x,A81x,A82x,A83x,A84x,A85x,A86x,A87x,A88x,A89x,A90x,A91x,A92x,A93x,A94x,A95x,A96x,A97x,A98x,A99x,A100x,A101x,A102x,A103x,A104x,A105x,A106x,A107x,A108x,A109x,A110x,A111x,A112x,A113x,A114x,A115x,A116x,A117x,A118x,A119x,A120x,A121x,A122x,A123x,A124x,A125x,A126x,A127x,A128x,A129x,A130x,A131x,A132x,A133x,A134x,A135x,A136x,A137x,A138x,A139x,A140x,A141x,A142x,A143x,A144x,A145x,A146x,A147x,A148x,A149x,A150x,A151x,A152x,A153x,A154x,A155x,A156x,A157x,A158x,A159x,A160x,A161x,A162x,A163x,A164x,A165x,A166x,A167x,A168x,A169x,A170x,A171x,A172x,A173x,A174x,A175x,A176x,A177x,A178x,A179x,A180x,A181x,A182x,A183x,A184x,A185x,A186x);
	input clk;
	input reset;
	input [7:0] A0x;
	input [7:0] A1x;
	input [7:0] A2x;
	input [7:0] A3x;
	input [7:0] A4x;
	input [7:0] A5x;
	input [7:0] A6x;
	input [7:0] A7x;
	input [7:0] A8x;
	input [7:0] A9x;
	input [7:0] A10x;
	input [7:0] A11x;
	input [7:0] A12x;
	input [7:0] A13x;
	input [7:0] A14x;
	input [7:0] A15x;
	input [7:0] A16x;
	input [7:0] A17x;
	input [7:0] A18x;
	input [7:0] A19x;
	input [7:0] A20x;
	input [7:0] A21x;
	input [7:0] A22x;
	input [7:0] A23x;
	input [7:0] A24x;
	input [7:0] A25x;
	input [7:0] A26x;
	input [7:0] A27x;
	input [7:0] A28x;
	input [7:0] A29x;
	input [7:0] A30x;
	input [7:0] A31x;
	input [7:0] A32x;
	input [7:0] A33x;
	input [7:0] A34x;
	input [7:0] A35x;
	input [7:0] A36x;
	input [7:0] A37x;
	input [7:0] A38x;
	input [7:0] A39x;
	input [7:0] A40x;
	input [7:0] A41x;
	input [7:0] A42x;
	input [7:0] A43x;
	input [7:0] A44x;
	input [7:0] A45x;
	input [7:0] A46x;
	input [7:0] A47x;
	input [7:0] A48x;
	input [7:0] A49x;
	input [7:0] A50x;
	input [7:0] A51x;
	input [7:0] A52x;
	input [7:0] A53x;
	input [7:0] A54x;
	input [7:0] A55x;
	input [7:0] A56x;
	input [7:0] A57x;
	input [7:0] A58x;
	input [7:0] A59x;
	input [7:0] A60x;
	input [7:0] A61x;
	input [7:0] A62x;
	input [7:0] A63x;
	input [7:0] A64x;
	input [7:0] A65x;
	input [7:0] A66x;
	input [7:0] A67x;
	input [7:0] A68x;
	input [7:0] A69x;
	input [7:0] A70x;
	input [7:0] A71x;
	input [7:0] A72x;
	input [7:0] A73x;
	input [7:0] A74x;
	input [7:0] A75x;
	input [7:0] A76x;
	input [7:0] A77x;
	input [7:0] A78x;
	input [7:0] A79x;
	input [7:0] A80x;
	input [7:0] A81x;
	input [7:0] A82x;
	input [7:0] A83x;
	input [7:0] A84x;
	input [7:0] A85x;
	input [7:0] A86x;
	input [7:0] A87x;
	input [7:0] A88x;
	input [7:0] A89x;
	input [7:0] A90x;
	input [7:0] A91x;
	input [7:0] A92x;
	input [7:0] A93x;
	input [7:0] A94x;
	input [7:0] A95x;
	input [7:0] A96x;
	input [7:0] A97x;
	input [7:0] A98x;
	input [7:0] A99x;
	input [7:0] A100x;
	input [7:0] A101x;
	input [7:0] A102x;
	input [7:0] A103x;
	input [7:0] A104x;
	input [7:0] A105x;
	input [7:0] A106x;
	input [7:0] A107x;
	input [7:0] A108x;
	input [7:0] A109x;
	input [7:0] A110x;
	input [7:0] A111x;
	input [7:0] A112x;
	input [7:0] A113x;
	input [7:0] A114x;
	input [7:0] A115x;
	input [7:0] A116x;
	input [7:0] A117x;
	input [7:0] A118x;
	input [7:0] A119x;
	input [7:0] A120x;
	input [7:0] A121x;
	input [7:0] A122x;
	input [7:0] A123x;
	input [7:0] A124x;
	input [7:0] A125x;
	input [7:0] A126x;
	input [7:0] A127x;
	input [7:0] A128x;
	input [7:0] A129x;
	input [7:0] A130x;
	input [7:0] A131x;
	input [7:0] A132x;
	input [7:0] A133x;
	input [7:0] A134x;
	input [7:0] A135x;
	input [7:0] A136x;
	input [7:0] A137x;
	input [7:0] A138x;
	input [7:0] A139x;
	input [7:0] A140x;
	input [7:0] A141x;
	input [7:0] A142x;
	input [7:0] A143x;
	input [7:0] A144x;
	input [7:0] A145x;
	input [7:0] A146x;
	input [7:0] A147x;
	input [7:0] A148x;
	input [7:0] A149x;
	input [7:0] A150x;
	input [7:0] A151x;
	input [7:0] A152x;
	input [7:0] A153x;
	input [7:0] A154x;
	input [7:0] A155x;
	input [7:0] A156x;
	input [7:0] A157x;
	input [7:0] A158x;
	input [7:0] A159x;
	input [7:0] A160x;
	input [7:0] A161x;
	input [7:0] A162x;
	input [7:0] A163x;
	input [7:0] A164x;
	input [7:0] A165x;
	input [7:0] A166x;
	input [7:0] A167x;
	input [7:0] A168x;
	input [7:0] A169x;
	input [7:0] A170x;
	input [7:0] A171x;
	input [7:0] A172x;
	input [7:0] A173x;
	input [7:0] A174x;
	input [7:0] A175x;
	input [7:0] A176x;
	input [7:0] A177x;
	input [7:0] A178x;
	input [7:0] A179x;
	input [7:0] A180x;
	input [7:0] A181x;
	input [7:0] A182x;
	input [7:0] A183x;
	input [7:0] A184x;
	input [7:0] A185x;
	input [7:0] A186x;
	reg signed [7:0] A0x_c;
	reg signed [7:0] A1x_c;
	reg signed [7:0] A2x_c;
	reg signed [7:0] A3x_c;
	reg signed [7:0] A4x_c;
	reg signed [7:0] A5x_c;
	reg signed [7:0] A6x_c;
	reg signed [7:0] A7x_c;
	reg signed [7:0] A8x_c;
	reg signed [7:0] A9x_c;
	reg signed [7:0] A10x_c;
	reg signed [7:0] A11x_c;
	reg signed [7:0] A12x_c;
	reg signed [7:0] A13x_c;
	reg signed [7:0] A14x_c;
	reg signed [7:0] A15x_c;
	reg signed [7:0] A16x_c;
	reg signed [7:0] A17x_c;
	reg signed [7:0] A18x_c;
	reg signed [7:0] A19x_c;
	reg signed [7:0] A20x_c;
	reg signed [7:0] A21x_c;
	reg signed [7:0] A22x_c;
	reg signed [7:0] A23x_c;
	reg signed [7:0] A24x_c;
	reg signed [7:0] A25x_c;
	reg signed [7:0] A26x_c;
	reg signed [7:0] A27x_c;
	reg signed [7:0] A28x_c;
	reg signed [7:0] A29x_c;
	reg signed [7:0] A30x_c;
	reg signed [7:0] A31x_c;
	reg signed [7:0] A32x_c;
	reg signed [7:0] A33x_c;
	reg signed [7:0] A34x_c;
	reg signed [7:0] A35x_c;
	reg signed [7:0] A36x_c;
	reg signed [7:0] A37x_c;
	reg signed [7:0] A38x_c;
	reg signed [7:0] A39x_c;
	reg signed [7:0] A40x_c;
	reg signed [7:0] A41x_c;
	reg signed [7:0] A42x_c;
	reg signed [7:0] A43x_c;
	reg signed [7:0] A44x_c;
	reg signed [7:0] A45x_c;
	reg signed [7:0] A46x_c;
	reg signed [7:0] A47x_c;
	reg signed [7:0] A48x_c;
	reg signed [7:0] A49x_c;
	reg signed [7:0] A50x_c;
	reg signed [7:0] A51x_c;
	reg signed [7:0] A52x_c;
	reg signed [7:0] A53x_c;
	reg signed [7:0] A54x_c;
	reg signed [7:0] A55x_c;
	reg signed [7:0] A56x_c;
	reg signed [7:0] A57x_c;
	reg signed [7:0] A58x_c;
	reg signed [7:0] A59x_c;
	reg signed [7:0] A60x_c;
	reg signed [7:0] A61x_c;
	reg signed [7:0] A62x_c;
	reg signed [7:0] A63x_c;
	reg signed [7:0] A64x_c;
	reg signed [7:0] A65x_c;
	reg signed [7:0] A66x_c;
	reg signed [7:0] A67x_c;
	reg signed [7:0] A68x_c;
	reg signed [7:0] A69x_c;
	reg signed [7:0] A70x_c;
	reg signed [7:0] A71x_c;
	reg signed [7:0] A72x_c;
	reg signed [7:0] A73x_c;
	reg signed [7:0] A74x_c;
	reg signed [7:0] A75x_c;
	reg signed [7:0] A76x_c;
	reg signed [7:0] A77x_c;
	reg signed [7:0] A78x_c;
	reg signed [7:0] A79x_c;
	reg signed [7:0] A80x_c;
	reg signed [7:0] A81x_c;
	reg signed [7:0] A82x_c;
	reg signed [7:0] A83x_c;
	reg signed [7:0] A84x_c;
	reg signed [7:0] A85x_c;
	reg signed [7:0] A86x_c;
	reg signed [7:0] A87x_c;
	reg signed [7:0] A88x_c;
	reg signed [7:0] A89x_c;
	reg signed [7:0] A90x_c;
	reg signed [7:0] A91x_c;
	reg signed [7:0] A92x_c;
	reg signed [7:0] A93x_c;
	reg signed [7:0] A94x_c;
	reg signed [7:0] A95x_c;
	reg signed [7:0] A96x_c;
	reg signed [7:0] A97x_c;
	reg signed [7:0] A98x_c;
	reg signed [7:0] A99x_c;
	reg signed [7:0] A100x_c;
	reg signed [7:0] A101x_c;
	reg signed [7:0] A102x_c;
	reg signed [7:0] A103x_c;
	reg signed [7:0] A104x_c;
	reg signed [7:0] A105x_c;
	reg signed [7:0] A106x_c;
	reg signed [7:0] A107x_c;
	reg signed [7:0] A108x_c;
	reg signed [7:0] A109x_c;
	reg signed [7:0] A110x_c;
	reg signed [7:0] A111x_c;
	reg signed [7:0] A112x_c;
	reg signed [7:0] A113x_c;
	reg signed [7:0] A114x_c;
	reg signed [7:0] A115x_c;
	reg signed [7:0] A116x_c;
	reg signed [7:0] A117x_c;
	reg signed [7:0] A118x_c;
	reg signed [7:0] A119x_c;
	reg signed [7:0] A120x_c;
	reg signed [7:0] A121x_c;
	reg signed [7:0] A122x_c;
	reg signed [7:0] A123x_c;
	reg signed [7:0] A124x_c;
	reg signed [7:0] A125x_c;
	reg signed [7:0] A126x_c;
	reg signed [7:0] A127x_c;
	reg signed [7:0] A128x_c;
	reg signed [7:0] A129x_c;
	reg signed [7:0] A130x_c;
	reg signed [7:0] A131x_c;
	reg signed [7:0] A132x_c;
	reg signed [7:0] A133x_c;
	reg signed [7:0] A134x_c;
	reg signed [7:0] A135x_c;
	reg signed [7:0] A136x_c;
	reg signed [7:0] A137x_c;
	reg signed [7:0] A138x_c;
	reg signed [7:0] A139x_c;
	reg signed [7:0] A140x_c;
	reg signed [7:0] A141x_c;
	reg signed [7:0] A142x_c;
	reg signed [7:0] A143x_c;
	reg signed [7:0] A144x_c;
	reg signed [7:0] A145x_c;
	reg signed [7:0] A146x_c;
	reg signed [7:0] A147x_c;
	reg signed [7:0] A148x_c;
	reg signed [7:0] A149x_c;
	reg signed [7:0] A150x_c;
	reg signed [7:0] A151x_c;
	reg signed [7:0] A152x_c;
	reg signed [7:0] A153x_c;
	reg signed [7:0] A154x_c;
	reg signed [7:0] A155x_c;
	reg signed [7:0] A156x_c;
	reg signed [7:0] A157x_c;
	reg signed [7:0] A158x_c;
	reg signed [7:0] A159x_c;
	reg signed [7:0] A160x_c;
	reg signed [7:0] A161x_c;
	reg signed [7:0] A162x_c;
	reg signed [7:0] A163x_c;
	reg signed [7:0] A164x_c;
	reg signed [7:0] A165x_c;
	reg signed [7:0] A166x_c;
	reg signed [7:0] A167x_c;
	reg signed [7:0] A168x_c;
	reg signed [7:0] A169x_c;
	reg signed [7:0] A170x_c;
	reg signed [7:0] A171x_c;
	reg signed [7:0] A172x_c;
	reg signed [7:0] A173x_c;
	reg signed [7:0] A174x_c;
	reg signed [7:0] A175x_c;
	reg signed [7:0] A176x_c;
	reg signed [7:0] A177x_c;
	reg signed [7:0] A178x_c;
	reg signed [7:0] A179x_c;
	reg signed [7:0] A180x_c;
	reg signed [7:0] A181x_c;
	reg signed [7:0] A182x_c;
	reg signed [7:0] A183x_c;
	reg signed [7:0] A184x_c;
	reg signed [7:0] A185x_c;
	reg signed [7:0] A186x_c;
	wire [15:0] sum0x;
	wire [15:0] sum1x;
	wire [15:0] sum2x;
	wire [15:0] sum3x;
	wire [15:0] sum4x;
	wire [15:0] sum5x;
	wire [15:0] sum6x;
	wire [15:0] sum7x;
	wire [15:0] sum8x;
	wire [15:0] sum9x;
	wire [15:0] sum10x;
	wire [15:0] sum11x;
	wire [15:0] sum12x;
	wire [15:0] sum13x;
	wire [15:0] sum14x;
	wire [15:0] sum15x;
	wire [15:0] sum16x;
	wire [15:0] sum17x;
	wire [15:0] sum18x;
	wire [15:0] sum19x;
	wire [15:0] sum20x;
	wire [15:0] sum21x;
	wire [15:0] sum22x;
	wire [15:0] sum23x;
	wire [15:0] sum24x;
	wire [15:0] sum25x;
	wire [15:0] sum26x;
	wire [15:0] sum27x;
	wire [15:0] sum28x;
	wire [15:0] sum29x;
	wire [15:0] sum30x;
	wire [15:0] sum31x;
	wire [15:0] sum32x;
	wire [15:0] sum33x;
	wire [15:0] sum34x;
	wire [15:0] sum35x;
	wire [15:0] sum36x;
	wire [15:0] sum37x;
	wire [15:0] sum38x;
	wire [15:0] sum39x;
	wire [15:0] sum40x;
	wire [15:0] sum41x;
	wire [15:0] sum42x;
	wire [15:0] sum43x;
	wire [15:0] sum44x;
	wire [15:0] sum45x;
	wire [15:0] sum46x;
	wire [15:0] sum47x;
	wire [15:0] sum48x;
	wire [15:0] sum49x;
	wire [15:0] sum50x;
	wire [15:0] sum51x;
	wire [15:0] sum52x;
	wire [15:0] sum53x;
	wire [15:0] sum54x;
	wire [15:0] sum55x;
	wire [15:0] sum56x;
	wire [15:0] sum57x;
	wire [15:0] sum58x;
	wire [15:0] sum59x;
	wire [15:0] sum60x;
	wire [15:0] sum61x;
	wire [15:0] sum62x;
	wire [15:0] sum63x;
	wire [15:0] sum64x;
	wire [15:0] sum65x;
	wire [15:0] sum66x;
	wire [15:0] sum67x;
	wire [15:0] sum68x;
	wire [15:0] sum69x;
	wire [15:0] sum70x;
	wire [15:0] sum71x;
	wire [15:0] sum72x;
	wire [15:0] sum73x;
	wire [15:0] sum74x;
	wire [15:0] sum75x;
	wire [15:0] sum76x;
	wire [15:0] sum77x;
	wire [15:0] sum78x;
	wire [15:0] sum79x;
	wire [15:0] sum80x;
	wire [15:0] sum81x;
	wire [15:0] sum82x;
	wire [15:0] sum83x;
	wire [15:0] sum84x;
	wire [15:0] sum85x;
	wire [15:0] sum86x;
	wire [15:0] sum87x;
	wire [15:0] sum88x;
	wire [15:0] sum89x;
	wire [15:0] sum90x;
	wire [15:0] sum91x;
	wire [15:0] sum92x;
	wire [15:0] sum93x;
	wire [15:0] sum94x;
	wire [15:0] sum95x;
	wire [15:0] sum96x;
	wire [15:0] sum97x;
	wire [15:0] sum98x;
	wire [15:0] sum99x;
	wire [15:0] sum100x;
	wire [15:0] sum101x;
	wire [15:0] sum102x;
	wire [15:0] sum103x;
	wire [15:0] sum104x;
	wire [15:0] sum105x;
	wire [15:0] sum106x;
	wire [15:0] sum107x;
	wire [15:0] sum108x;
	wire [15:0] sum109x;
	wire [15:0] sum110x;
	wire [15:0] sum111x;
	wire [15:0] sum112x;
	wire [15:0] sum113x;
	wire [15:0] sum114x;
	wire [15:0] sum115x;
	wire [15:0] sum116x;
	wire [15:0] sum117x;
	wire [15:0] sum118x;
	wire [15:0] sum119x;
	wire [15:0] sum120x;
	wire [15:0] sum121x;
	wire [15:0] sum122x;
	wire [15:0] sum123x;
	wire [15:0] sum124x;
	wire [15:0] sum125x;
	wire [15:0] sum126x;
	wire [15:0] sum127x;
	wire [15:0] sum128x;
	wire [15:0] sum129x;
	wire [15:0] sum130x;
	wire [15:0] sum131x;
	wire [15:0] sum132x;
	wire [15:0] sum133x;
	wire [15:0] sum134x;
	wire [15:0] sum135x;
	wire [15:0] sum136x;
	wire [15:0] sum137x;
	wire [15:0] sum138x;
	wire [15:0] sum139x;
	wire [15:0] sum140x;
	wire [15:0] sum141x;
	wire [15:0] sum142x;
	wire [15:0] sum143x;
	wire [15:0] sum144x;
	wire [15:0] sum145x;
	wire [15:0] sum146x;
	wire [15:0] sum147x;
	wire [15:0] sum148x;
	wire [15:0] sum149x;
	wire [15:0] sum150x;
	wire [15:0] sum151x;
	wire [15:0] sum152x;
	wire [15:0] sum153x;
	wire [15:0] sum154x;
	wire [15:0] sum155x;
	wire [15:0] sum156x;
	wire [15:0] sum157x;
	wire [15:0] sum158x;
	wire [15:0] sum159x;
	wire [15:0] sum160x;
	wire [15:0] sum161x;
	wire [15:0] sum162x;
	wire [15:0] sum163x;
	wire [15:0] sum164x;
	wire [15:0] sum165x;
	wire [15:0] sum166x;
	wire [15:0] sum167x;
	wire [15:0] sum168x;
	wire [15:0] sum169x;
	wire [15:0] sum170x;
	wire [15:0] sum171x;
	wire [15:0] sum172x;
	wire [15:0] sum173x;
	wire [15:0] sum174x;
	wire [15:0] sum175x;
	wire [15:0] sum176x;
	wire [15:0] sum177x;
	wire [15:0] sum178x;
	wire [15:0] sum179x;
	wire [15:0] sum180x;
	wire [15:0] sum181x;
	wire [15:0] sum182x;
	wire [15:0] sum183x;
	wire [15:0] sum184x;
	wire [15:0] sum185x;
	wire [15:0] sum186x;
	output reg [7:0] N1x;
	reg signed [22:0] sumout;

	parameter signed [7:0] W0x=-8'd4;
	parameter signed [7:0] W1x=8'd38;
	parameter signed [7:0] W2x=-8'd40;
	parameter signed [7:0] W3x=-8'd36;
	parameter signed [7:0] W4x=-8'd62;
	parameter signed [7:0] W5x=-8'd18;
	parameter signed [7:0] W6x=8'd20;
	parameter signed [7:0] W7x=8'd20;
	parameter signed [7:0] W8x=8'd14;
	parameter signed [7:0] W9x=8'd18;
	parameter signed [7:0] W10x=-8'd2;
	parameter signed [7:0] W11x=8'd12;
	parameter signed [7:0] W12x=-8'd2;
	parameter signed [7:0] W13x=-8'd4;
	parameter signed [7:0] W14x=-8'd4;
	parameter signed [7:0] W15x=8'd4;
	parameter signed [7:0] W16x=-8'd4;
	parameter signed [7:0] W17x=8'd8;
	parameter signed [7:0] W18x=-8'd2;
	parameter signed [7:0] W19x=8'd2;
	parameter signed [7:0] W20x=-8'd2;
	parameter signed [7:0] W21x=-8'd4;
	parameter signed [7:0] W22x=-8'd6;
	parameter signed [7:0] W23x=-8'd6;
	parameter signed [7:0] W24x=8'd2;
	parameter signed [7:0] W25x=-8'd4;
	parameter signed [7:0] W26x=8'd2;
	parameter signed [7:0] W27x=8'd4;
	parameter signed [7:0] W28x=8'd8;
	parameter signed [7:0] W29x=8'd4;
	parameter signed [7:0] W30x=8'd6;
	parameter signed [7:0] W31x=8'd8;
	parameter signed [7:0] W32x=8'd4;
	parameter signed [7:0] W33x=-8'd4;
	parameter signed [7:0] W34x=-8'd4;
	parameter signed [7:0] W35x=-8'd16;
	parameter signed [7:0] W36x=-8'd6;
	parameter signed [7:0] W37x=8'd4;
	parameter signed [7:0] W38x=8'd2;
	parameter signed [7:0] W39x=8'd10;
	parameter signed [7:0] W40x=8'd12;
	parameter signed [7:0] W41x=8'd6;
	parameter signed [7:0] W42x=8'd8;
	parameter signed [7:0] W43x=8'd2;
	parameter signed [7:0] W44x=-8'd10;
	parameter signed [7:0] W45x=-8'd2;
	parameter signed [7:0] W46x=8'd6;
	parameter signed [7:0] W47x=-8'd24;
	parameter signed [7:0] W48x=-8'd22;
	parameter signed [7:0] W49x=-8'd8;
	parameter signed [7:0] W50x=-8'd12;
	parameter signed [7:0] W51x=-8'd16;
	parameter signed [7:0] W52x=-8'd14;
	parameter signed [7:0] W53x=-8'd12;
	parameter signed [7:0] W54x=-8'd8;
	parameter signed [7:0] W55x=8'd0;
	parameter signed [7:0] W56x=8'd2;
	parameter signed [7:0] W57x=-8'd2;
	parameter signed [7:0] W58x=8'd0;
	parameter signed [7:0] W59x=8'd6;
	parameter signed [7:0] W60x=8'd8;
	parameter signed [7:0] W61x=8'd6;
	parameter signed [7:0] W62x=8'd0;
	parameter signed [7:0] W63x=8'd4;
	parameter signed [7:0] W64x=8'd0;
	parameter signed [7:0] W65x=8'd10;
	parameter signed [7:0] W66x=8'd6;
	parameter signed [7:0] W67x=-8'd2;
	parameter signed [7:0] W68x=-8'd6;
	parameter signed [7:0] W69x=-8'd18;
	parameter signed [7:0] W70x=-8'd2;
	parameter signed [7:0] W71x=-8'd14;
	parameter signed [7:0] W72x=-8'd2;
	parameter signed [7:0] W73x=8'd10;
	parameter signed [7:0] W74x=8'd8;
	parameter signed [7:0] W75x=8'd14;
	parameter signed [7:0] W76x=8'd6;
	parameter signed [7:0] W77x=8'd12;
	parameter signed [7:0] W78x=8'd8;
	parameter signed [7:0] W79x=8'd10;
	parameter signed [7:0] W80x=8'd4;
	parameter signed [7:0] W81x=8'd0;
	parameter signed [7:0] W82x=8'd2;
	parameter signed [7:0] W83x=-8'd8;
	parameter signed [7:0] W84x=-8'd14;
	parameter signed [7:0] W85x=-8'd2;
	parameter signed [7:0] W86x=-8'd6;
	parameter signed [7:0] W87x=8'd12;
	parameter signed [7:0] W88x=-8'd4;
	parameter signed [7:0] W89x=8'd0;
	parameter signed [7:0] W90x=8'd6;
	parameter signed [7:0] W91x=-8'd2;
	parameter signed [7:0] W92x=8'd0;
	parameter signed [7:0] W93x=8'd4;
	parameter signed [7:0] W94x=-8'd4;
	parameter signed [7:0] W95x=-8'd14;
	parameter signed [7:0] W96x=-8'd4;
	parameter signed [7:0] W97x=-8'd14;
	parameter signed [7:0] W98x=-8'd6;
	parameter signed [7:0] W99x=-8'd4;
	parameter signed [7:0] W100x=8'd4;
	parameter signed [7:0] W101x=-8'd10;
	parameter signed [7:0] W102x=8'd0;
	parameter signed [7:0] W103x=8'd2;
	parameter signed [7:0] W104x=-8'd8;
	parameter signed [7:0] W105x=-8'd2;
	parameter signed [7:0] W106x=8'd4;
	parameter signed [7:0] W107x=8'd8;
	parameter signed [7:0] W108x=-8'd2;
	parameter signed [7:0] W109x=8'd2;
	parameter signed [7:0] W110x=8'd2;
	parameter signed [7:0] W111x=8'd6;
	parameter signed [7:0] W112x=8'd10;
	parameter signed [7:0] W113x=8'd0;
	parameter signed [7:0] W114x=8'd12;
	parameter signed [7:0] W115x=8'd4;
	parameter signed [7:0] W116x=8'd4;
	parameter signed [7:0] W117x=8'd4;
	parameter signed [7:0] W118x=8'd8;
	parameter signed [7:0] W119x=8'd2;
	parameter signed [7:0] W120x=8'd6;
	parameter signed [7:0] W121x=8'd4;
	parameter signed [7:0] W122x=8'd6;
	parameter signed [7:0] W123x=8'd0;
	parameter signed [7:0] W124x=8'd6;
	parameter signed [7:0] W125x=8'd6;
	parameter signed [7:0] W126x=8'd4;
	parameter signed [7:0] W127x=8'd4;
	parameter signed [7:0] W128x=8'd4;
	parameter signed [7:0] W129x=-8'd6;
	parameter signed [7:0] W130x=8'd2;
	parameter signed [7:0] W131x=8'd12;
	parameter signed [7:0] W132x=8'd0;
	parameter signed [7:0] W133x=8'd2;
	parameter signed [7:0] W134x=8'd6;
	parameter signed [7:0] W135x=8'd0;
	parameter signed [7:0] W136x=8'd6;
	parameter signed [7:0] W137x=8'd2;
	parameter signed [7:0] W138x=8'd6;
	parameter signed [7:0] W139x=8'd16;
	parameter signed [7:0] W140x=8'd4;
	parameter signed [7:0] W141x=8'd0;
	parameter signed [7:0] W142x=8'd0;
	parameter signed [7:0] W143x=8'd18;
	parameter signed [7:0] W144x=-8'd4;
	parameter signed [7:0] W145x=8'd4;
	parameter signed [7:0] W146x=8'd18;
	parameter signed [7:0] W147x=8'd6;
	parameter signed [7:0] W148x=8'd8;
	parameter signed [7:0] W149x=-8'd2;
	parameter signed [7:0] W150x=8'd18;
	parameter signed [7:0] W151x=-8'd6;
	parameter signed [7:0] W152x=8'd12;
	parameter signed [7:0] W153x=-8'd4;
	parameter signed [7:0] W154x=8'd12;
	parameter signed [7:0] W155x=8'd8;
	parameter signed [7:0] W156x=-8'd2;
	parameter signed [7:0] W157x=8'd2;
	parameter signed [7:0] W158x=8'd22;
	parameter signed [7:0] W159x=-8'd4;
	parameter signed [7:0] W160x=8'd4;
	parameter signed [7:0] W161x=-8'd2;
	parameter signed [7:0] W162x=-8'd18;
	parameter signed [7:0] W163x=8'd6;
	parameter signed [7:0] W164x=-8'd10;
	parameter signed [7:0] W165x=-8'd36;
	parameter signed [7:0] W166x=-8'd36;
	parameter signed [7:0] W167x=-8'd4;
	parameter signed [7:0] W168x=-8'd4;
	parameter signed [7:0] W169x=-8'd18;
	parameter signed [7:0] W170x=-8'd20;
	parameter signed [7:0] W171x=-8'd10;
	parameter signed [7:0] W172x=-8'd38;
	parameter signed [7:0] W173x=8'd38;
	parameter signed [7:0] W174x=8'd18;
	parameter signed [7:0] W175x=8'd40;
	parameter signed [7:0] W176x=8'd20;
	parameter signed [7:0] W177x=8'd42;
	parameter signed [7:0] W178x=8'd24;
	parameter signed [7:0] W179x=8'd6;
	parameter signed [7:0] W180x=8'd8;
	parameter signed [7:0] W181x=8'd0;
	parameter signed [7:0] W182x=-8'd4;
	parameter signed [7:0] W183x=8'd44;
	parameter signed [7:0] W184x=8'd62;
	parameter signed [7:0] W185x=8'd62;
	parameter signed [7:0] W186x=8'd4;
	parameter [15:0] B0x=16'd0;


	assign sum0x = A0x_c*W0x;
	assign sum1x = A1x_c*W1x;
	assign sum2x = A2x_c*W2x;
	assign sum3x = A3x_c*W3x;
	assign sum4x = A4x_c*W4x;
	assign sum5x = A5x_c*W5x;
	assign sum6x = A6x_c*W6x;
	assign sum7x = A7x_c*W7x;
	assign sum8x = A8x_c*W8x;
	assign sum9x = A9x_c*W9x;
	assign sum10x = A10x_c*W10x;
	assign sum11x = A11x_c*W11x;
	assign sum12x = A12x_c*W12x;
	assign sum13x = A13x_c*W13x;
	assign sum14x = A14x_c*W14x;
	assign sum15x = A15x_c*W15x;
	assign sum16x = A16x_c*W16x;
	assign sum17x = A17x_c*W17x;
	assign sum18x = A18x_c*W18x;
	assign sum19x = A19x_c*W19x;
	assign sum20x = A20x_c*W20x;
	assign sum21x = A21x_c*W21x;
	assign sum22x = A22x_c*W22x;
	assign sum23x = A23x_c*W23x;
	assign sum24x = A24x_c*W24x;
	assign sum25x = A25x_c*W25x;
	assign sum26x = A26x_c*W26x;
	assign sum27x = A27x_c*W27x;
	assign sum28x = A28x_c*W28x;
	assign sum29x = A29x_c*W29x;
	assign sum30x = A30x_c*W30x;
	assign sum31x = A31x_c*W31x;
	assign sum32x = A32x_c*W32x;
	assign sum33x = A33x_c*W33x;
	assign sum34x = A34x_c*W34x;
	assign sum35x = A35x_c*W35x;
	assign sum36x = A36x_c*W36x;
	assign sum37x = A37x_c*W37x;
	assign sum38x = A38x_c*W38x;
	assign sum39x = A39x_c*W39x;
	assign sum40x = A40x_c*W40x;
	assign sum41x = A41x_c*W41x;
	assign sum42x = A42x_c*W42x;
	assign sum43x = A43x_c*W43x;
	assign sum44x = A44x_c*W44x;
	assign sum45x = A45x_c*W45x;
	assign sum46x = A46x_c*W46x;
	assign sum47x = A47x_c*W47x;
	assign sum48x = A48x_c*W48x;
	assign sum49x = A49x_c*W49x;
	assign sum50x = A50x_c*W50x;
	assign sum51x = A51x_c*W51x;
	assign sum52x = A52x_c*W52x;
	assign sum53x = A53x_c*W53x;
	assign sum54x = A54x_c*W54x;
	assign sum55x = A55x_c*W55x;
	assign sum56x = A56x_c*W56x;
	assign sum57x = A57x_c*W57x;
	assign sum58x = A58x_c*W58x;
	assign sum59x = A59x_c*W59x;
	assign sum60x = A60x_c*W60x;
	assign sum61x = A61x_c*W61x;
	assign sum62x = A62x_c*W62x;
	assign sum63x = A63x_c*W63x;
	assign sum64x = A64x_c*W64x;
	assign sum65x = A65x_c*W65x;
	assign sum66x = A66x_c*W66x;
	assign sum67x = A67x_c*W67x;
	assign sum68x = A68x_c*W68x;
	assign sum69x = A69x_c*W69x;
	assign sum70x = A70x_c*W70x;
	assign sum71x = A71x_c*W71x;
	assign sum72x = A72x_c*W72x;
	assign sum73x = A73x_c*W73x;
	assign sum74x = A74x_c*W74x;
	assign sum75x = A75x_c*W75x;
	assign sum76x = A76x_c*W76x;
	assign sum77x = A77x_c*W77x;
	assign sum78x = A78x_c*W78x;
	assign sum79x = A79x_c*W79x;
	assign sum80x = A80x_c*W80x;
	assign sum81x = A81x_c*W81x;
	assign sum82x = A82x_c*W82x;
	assign sum83x = A83x_c*W83x;
	assign sum84x = A84x_c*W84x;
	assign sum85x = A85x_c*W85x;
	assign sum86x = A86x_c*W86x;
	assign sum87x = A87x_c*W87x;
	assign sum88x = A88x_c*W88x;
	assign sum89x = A89x_c*W89x;
	assign sum90x = A90x_c*W90x;
	assign sum91x = A91x_c*W91x;
	assign sum92x = A92x_c*W92x;
	assign sum93x = A93x_c*W93x;
	assign sum94x = A94x_c*W94x;
	assign sum95x = A95x_c*W95x;
	assign sum96x = A96x_c*W96x;
	assign sum97x = A97x_c*W97x;
	assign sum98x = A98x_c*W98x;
	assign sum99x = A99x_c*W99x;
	assign sum100x = A100x_c*W100x;
	assign sum101x = A101x_c*W101x;
	assign sum102x = A102x_c*W102x;
	assign sum103x = A103x_c*W103x;
	assign sum104x = A104x_c*W104x;
	assign sum105x = A105x_c*W105x;
	assign sum106x = A106x_c*W106x;
	assign sum107x = A107x_c*W107x;
	assign sum108x = A108x_c*W108x;
	assign sum109x = A109x_c*W109x;
	assign sum110x = A110x_c*W110x;
	assign sum111x = A111x_c*W111x;
	assign sum112x = A112x_c*W112x;
	assign sum113x = A113x_c*W113x;
	assign sum114x = A114x_c*W114x;
	assign sum115x = A115x_c*W115x;
	assign sum116x = A116x_c*W116x;
	assign sum117x = A117x_c*W117x;
	assign sum118x = A118x_c*W118x;
	assign sum119x = A119x_c*W119x;
	assign sum120x = A120x_c*W120x;
	assign sum121x = A121x_c*W121x;
	assign sum122x = A122x_c*W122x;
	assign sum123x = A123x_c*W123x;
	assign sum124x = A124x_c*W124x;
	assign sum125x = A125x_c*W125x;
	assign sum126x = A126x_c*W126x;
	assign sum127x = A127x_c*W127x;
	assign sum128x = A128x_c*W128x;
	assign sum129x = A129x_c*W129x;
	assign sum130x = A130x_c*W130x;
	assign sum131x = A131x_c*W131x;
	assign sum132x = A132x_c*W132x;
	assign sum133x = A133x_c*W133x;
	assign sum134x = A134x_c*W134x;
	assign sum135x = A135x_c*W135x;
	assign sum136x = A136x_c*W136x;
	assign sum137x = A137x_c*W137x;
	assign sum138x = A138x_c*W138x;
	assign sum139x = A139x_c*W139x;
	assign sum140x = A140x_c*W140x;
	assign sum141x = A141x_c*W141x;
	assign sum142x = A142x_c*W142x;
	assign sum143x = A143x_c*W143x;
	assign sum144x = A144x_c*W144x;
	assign sum145x = A145x_c*W145x;
	assign sum146x = A146x_c*W146x;
	assign sum147x = A147x_c*W147x;
	assign sum148x = A148x_c*W148x;
	assign sum149x = A149x_c*W149x;
	assign sum150x = A150x_c*W150x;
	assign sum151x = A151x_c*W151x;
	assign sum152x = A152x_c*W152x;
	assign sum153x = A153x_c*W153x;
	assign sum154x = A154x_c*W154x;
	assign sum155x = A155x_c*W155x;
	assign sum156x = A156x_c*W156x;
	assign sum157x = A157x_c*W157x;
	assign sum158x = A158x_c*W158x;
	assign sum159x = A159x_c*W159x;
	assign sum160x = A160x_c*W160x;
	assign sum161x = A161x_c*W161x;
	assign sum162x = A162x_c*W162x;
	assign sum163x = A163x_c*W163x;
	assign sum164x = A164x_c*W164x;
	assign sum165x = A165x_c*W165x;
	assign sum166x = A166x_c*W166x;
	assign sum167x = A167x_c*W167x;
	assign sum168x = A168x_c*W168x;
	assign sum169x = A169x_c*W169x;
	assign sum170x = A170x_c*W170x;
	assign sum171x = A171x_c*W171x;
	assign sum172x = A172x_c*W172x;
	assign sum173x = A173x_c*W173x;
	assign sum174x = A174x_c*W174x;
	assign sum175x = A175x_c*W175x;
	assign sum176x = A176x_c*W176x;
	assign sum177x = A177x_c*W177x;
	assign sum178x = A178x_c*W178x;
	assign sum179x = A179x_c*W179x;
	assign sum180x = A180x_c*W180x;
	assign sum181x = A181x_c*W181x;
	assign sum182x = A182x_c*W182x;
	assign sum183x = A183x_c*W183x;
	assign sum184x = A184x_c*W184x;
	assign sum185x = A185x_c*W185x;
	assign sum186x = A186x_c*W186x;

	always@(posedge clk) begin

		if(reset)
			begin
			N1x<=8'd0;
			sumout<=16'd0;
			A0x_c <= 8'd0;
			A1x_c <= 8'd0;
			A2x_c <= 8'd0;
			A3x_c <= 8'd0;
			A4x_c <= 8'd0;
			A5x_c <= 8'd0;
			A6x_c <= 8'd0;
			A7x_c <= 8'd0;
			A8x_c <= 8'd0;
			A9x_c <= 8'd0;
			A10x_c <= 8'd0;
			A11x_c <= 8'd0;
			A12x_c <= 8'd0;
			A13x_c <= 8'd0;
			A14x_c <= 8'd0;
			A15x_c <= 8'd0;
			A16x_c <= 8'd0;
			A17x_c <= 8'd0;
			A18x_c <= 8'd0;
			A19x_c <= 8'd0;
			A20x_c <= 8'd0;
			A21x_c <= 8'd0;
			A22x_c <= 8'd0;
			A23x_c <= 8'd0;
			A24x_c <= 8'd0;
			A25x_c <= 8'd0;
			A26x_c <= 8'd0;
			A27x_c <= 8'd0;
			A28x_c <= 8'd0;
			A29x_c <= 8'd0;
			A30x_c <= 8'd0;
			A31x_c <= 8'd0;
			A32x_c <= 8'd0;
			A33x_c <= 8'd0;
			A34x_c <= 8'd0;
			A35x_c <= 8'd0;
			A36x_c <= 8'd0;
			A37x_c <= 8'd0;
			A38x_c <= 8'd0;
			A39x_c <= 8'd0;
			A40x_c <= 8'd0;
			A41x_c <= 8'd0;
			A42x_c <= 8'd0;
			A43x_c <= 8'd0;
			A44x_c <= 8'd0;
			A45x_c <= 8'd0;
			A46x_c <= 8'd0;
			A47x_c <= 8'd0;
			A48x_c <= 8'd0;
			A49x_c <= 8'd0;
			A50x_c <= 8'd0;
			A51x_c <= 8'd0;
			A52x_c <= 8'd0;
			A53x_c <= 8'd0;
			A54x_c <= 8'd0;
			A55x_c <= 8'd0;
			A56x_c <= 8'd0;
			A57x_c <= 8'd0;
			A58x_c <= 8'd0;
			A59x_c <= 8'd0;
			A60x_c <= 8'd0;
			A61x_c <= 8'd0;
			A62x_c <= 8'd0;
			A63x_c <= 8'd0;
			A64x_c <= 8'd0;
			A65x_c <= 8'd0;
			A66x_c <= 8'd0;
			A67x_c <= 8'd0;
			A68x_c <= 8'd0;
			A69x_c <= 8'd0;
			A70x_c <= 8'd0;
			A71x_c <= 8'd0;
			A72x_c <= 8'd0;
			A73x_c <= 8'd0;
			A74x_c <= 8'd0;
			A75x_c <= 8'd0;
			A76x_c <= 8'd0;
			A77x_c <= 8'd0;
			A78x_c <= 8'd0;
			A79x_c <= 8'd0;
			A80x_c <= 8'd0;
			A81x_c <= 8'd0;
			A82x_c <= 8'd0;
			A83x_c <= 8'd0;
			A84x_c <= 8'd0;
			A85x_c <= 8'd0;
			A86x_c <= 8'd0;
			A87x_c <= 8'd0;
			A88x_c <= 8'd0;
			A89x_c <= 8'd0;
			A90x_c <= 8'd0;
			A91x_c <= 8'd0;
			A92x_c <= 8'd0;
			A93x_c <= 8'd0;
			A94x_c <= 8'd0;
			A95x_c <= 8'd0;
			A96x_c <= 8'd0;
			A97x_c <= 8'd0;
			A98x_c <= 8'd0;
			A99x_c <= 8'd0;
			A100x_c <= 8'd0;
			A101x_c <= 8'd0;
			A102x_c <= 8'd0;
			A103x_c <= 8'd0;
			A104x_c <= 8'd0;
			A105x_c <= 8'd0;
			A106x_c <= 8'd0;
			A107x_c <= 8'd0;
			A108x_c <= 8'd0;
			A109x_c <= 8'd0;
			A110x_c <= 8'd0;
			A111x_c <= 8'd0;
			A112x_c <= 8'd0;
			A113x_c <= 8'd0;
			A114x_c <= 8'd0;
			A115x_c <= 8'd0;
			A116x_c <= 8'd0;
			A117x_c <= 8'd0;
			A118x_c <= 8'd0;
			A119x_c <= 8'd0;
			A120x_c <= 8'd0;
			A121x_c <= 8'd0;
			A122x_c <= 8'd0;
			A123x_c <= 8'd0;
			A124x_c <= 8'd0;
			A125x_c <= 8'd0;
			A126x_c <= 8'd0;
			A127x_c <= 8'd0;
			A128x_c <= 8'd0;
			A129x_c <= 8'd0;
			A130x_c <= 8'd0;
			A131x_c <= 8'd0;
			A132x_c <= 8'd0;
			A133x_c <= 8'd0;
			A134x_c <= 8'd0;
			A135x_c <= 8'd0;
			A136x_c <= 8'd0;
			A137x_c <= 8'd0;
			A138x_c <= 8'd0;
			A139x_c <= 8'd0;
			A140x_c <= 8'd0;
			A141x_c <= 8'd0;
			A142x_c <= 8'd0;
			A143x_c <= 8'd0;
			A144x_c <= 8'd0;
			A145x_c <= 8'd0;
			A146x_c <= 8'd0;
			A147x_c <= 8'd0;
			A148x_c <= 8'd0;
			A149x_c <= 8'd0;
			A150x_c <= 8'd0;
			A151x_c <= 8'd0;
			A152x_c <= 8'd0;
			A153x_c <= 8'd0;
			A154x_c <= 8'd0;
			A155x_c <= 8'd0;
			A156x_c <= 8'd0;
			A157x_c <= 8'd0;
			A158x_c <= 8'd0;
			A159x_c <= 8'd0;
			A160x_c <= 8'd0;
			A161x_c <= 8'd0;
			A162x_c <= 8'd0;
			A163x_c <= 8'd0;
			A164x_c <= 8'd0;
			A165x_c <= 8'd0;
			A166x_c <= 8'd0;
			A167x_c <= 8'd0;
			A168x_c <= 8'd0;
			A169x_c <= 8'd0;
			A170x_c <= 8'd0;
			A171x_c <= 8'd0;
			A172x_c <= 8'd0;
			A173x_c <= 8'd0;
			A174x_c <= 8'd0;
			A175x_c <= 8'd0;
			A176x_c <= 8'd0;
			A177x_c <= 8'd0;
			A178x_c <= 8'd0;
			A179x_c <= 8'd0;
			A180x_c <= 8'd0;
			A181x_c <= 8'd0;
			A182x_c <= 8'd0;
			A183x_c <= 8'd0;
			A184x_c <= 8'd0;
			A185x_c <= 8'd0;
			A186x_c <= 8'd0;
			end
		else
			begin
			A0x_c <= A0x;
			A1x_c <= A1x;
			A2x_c <= A2x;
			A3x_c <= A3x;
			A4x_c <= A4x;
			A5x_c <= A5x;
			A6x_c <= A6x;
			A7x_c <= A7x;
			A8x_c <= A8x;
			A9x_c <= A9x;
			A10x_c <= A10x;
			A11x_c <= A11x;
			A12x_c <= A12x;
			A13x_c <= A13x;
			A14x_c <= A14x;
			A15x_c <= A15x;
			A16x_c <= A16x;
			A17x_c <= A17x;
			A18x_c <= A18x;
			A19x_c <= A19x;
			A20x_c <= A20x;
			A21x_c <= A21x;
			A22x_c <= A22x;
			A23x_c <= A23x;
			A24x_c <= A24x;
			A25x_c <= A25x;
			A26x_c <= A26x;
			A27x_c <= A27x;
			A28x_c <= A28x;
			A29x_c <= A29x;
			A30x_c <= A30x;
			A31x_c <= A31x;
			A32x_c <= A32x;
			A33x_c <= A33x;
			A34x_c <= A34x;
			A35x_c <= A35x;
			A36x_c <= A36x;
			A37x_c <= A37x;
			A38x_c <= A38x;
			A39x_c <= A39x;
			A40x_c <= A40x;
			A41x_c <= A41x;
			A42x_c <= A42x;
			A43x_c <= A43x;
			A44x_c <= A44x;
			A45x_c <= A45x;
			A46x_c <= A46x;
			A47x_c <= A47x;
			A48x_c <= A48x;
			A49x_c <= A49x;
			A50x_c <= A50x;
			A51x_c <= A51x;
			A52x_c <= A52x;
			A53x_c <= A53x;
			A54x_c <= A54x;
			A55x_c <= A55x;
			A56x_c <= A56x;
			A57x_c <= A57x;
			A58x_c <= A58x;
			A59x_c <= A59x;
			A60x_c <= A60x;
			A61x_c <= A61x;
			A62x_c <= A62x;
			A63x_c <= A63x;
			A64x_c <= A64x;
			A65x_c <= A65x;
			A66x_c <= A66x;
			A67x_c <= A67x;
			A68x_c <= A68x;
			A69x_c <= A69x;
			A70x_c <= A70x;
			A71x_c <= A71x;
			A72x_c <= A72x;
			A73x_c <= A73x;
			A74x_c <= A74x;
			A75x_c <= A75x;
			A76x_c <= A76x;
			A77x_c <= A77x;
			A78x_c <= A78x;
			A79x_c <= A79x;
			A80x_c <= A80x;
			A81x_c <= A81x;
			A82x_c <= A82x;
			A83x_c <= A83x;
			A84x_c <= A84x;
			A85x_c <= A85x;
			A86x_c <= A86x;
			A87x_c <= A87x;
			A88x_c <= A88x;
			A89x_c <= A89x;
			A90x_c <= A90x;
			A91x_c <= A91x;
			A92x_c <= A92x;
			A93x_c <= A93x;
			A94x_c <= A94x;
			A95x_c <= A95x;
			A96x_c <= A96x;
			A97x_c <= A97x;
			A98x_c <= A98x;
			A99x_c <= A99x;
			A100x_c <= A100x;
			A101x_c <= A101x;
			A102x_c <= A102x;
			A103x_c <= A103x;
			A104x_c <= A104x;
			A105x_c <= A105x;
			A106x_c <= A106x;
			A107x_c <= A107x;
			A108x_c <= A108x;
			A109x_c <= A109x;
			A110x_c <= A110x;
			A111x_c <= A111x;
			A112x_c <= A112x;
			A113x_c <= A113x;
			A114x_c <= A114x;
			A115x_c <= A115x;
			A116x_c <= A116x;
			A117x_c <= A117x;
			A118x_c <= A118x;
			A119x_c <= A119x;
			A120x_c <= A120x;
			A121x_c <= A121x;
			A122x_c <= A122x;
			A123x_c <= A123x;
			A124x_c <= A124x;
			A125x_c <= A125x;
			A126x_c <= A126x;
			A127x_c <= A127x;
			A128x_c <= A128x;
			A129x_c <= A129x;
			A130x_c <= A130x;
			A131x_c <= A131x;
			A132x_c <= A132x;
			A133x_c <= A133x;
			A134x_c <= A134x;
			A135x_c <= A135x;
			A136x_c <= A136x;
			A137x_c <= A137x;
			A138x_c <= A138x;
			A139x_c <= A139x;
			A140x_c <= A140x;
			A141x_c <= A141x;
			A142x_c <= A142x;
			A143x_c <= A143x;
			A144x_c <= A144x;
			A145x_c <= A145x;
			A146x_c <= A146x;
			A147x_c <= A147x;
			A148x_c <= A148x;
			A149x_c <= A149x;
			A150x_c <= A150x;
			A151x_c <= A151x;
			A152x_c <= A152x;
			A153x_c <= A153x;
			A154x_c <= A154x;
			A155x_c <= A155x;
			A156x_c <= A156x;
			A157x_c <= A157x;
			A158x_c <= A158x;
			A159x_c <= A159x;
			A160x_c <= A160x;
			A161x_c <= A161x;
			A162x_c <= A162x;
			A163x_c <= A163x;
			A164x_c <= A164x;
			A165x_c <= A165x;
			A166x_c <= A166x;
			A167x_c <= A167x;
			A168x_c <= A168x;
			A169x_c <= A169x;
			A170x_c <= A170x;
			A171x_c <= A171x;
			A172x_c <= A172x;
			A173x_c <= A173x;
			A174x_c <= A174x;
			A175x_c <= A175x;
			A176x_c <= A176x;
			A177x_c <= A177x;
			A178x_c <= A178x;
			A179x_c <= A179x;
			A180x_c <= A180x;
			A181x_c <= A181x;
			A182x_c <= A182x;
			A183x_c <= A183x;
			A184x_c <= A184x;
			A185x_c <= A185x;
			A186x_c <= A186x;
			sumout<={sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x}+{sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x}+{sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x}+{sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x}+{sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x}+{sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x}+{sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x}+{sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x}+{sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x}+{sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x}+{sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x}+{sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x}+{sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x}+{sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x}+{sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x}+{sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x}+{sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x}+{sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x}+{sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x}+{sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x}+{sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x}+{sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x}+{sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x}+{sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x}+{sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x}+{sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x}+{sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x}+{sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x}+{sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x}+{sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x}+{sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x}+{sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x}+{sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x}+{sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x}+{sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x}+{sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x}+{sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x}+{sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x}+{sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x}+{sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x}+{sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x}+{sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x}+{sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x}+{sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x}+{sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x}+{sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x}+{sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x}+{sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x}+{sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x}+{sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x}+{sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x}+{sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x}+{sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x}+{sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x}+{sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x}+{sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x}+{sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x}+{sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x}+{sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x}+{sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x}+{sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x}+{sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x}+{sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x}+{sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x}+{sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x}+{sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x}+{sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x}+{sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x}+{sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x}+{sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x}+{sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x}+{sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x}+{sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x}+{sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x}+{sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x}+{sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x}+{sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x}+{sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x}+{sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x}+{sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x}+{sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x}+{sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x}+{sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x}+{sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x}+{sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x}+{sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x}+{sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x}+{sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x}+{sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x}+{sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x}+{sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x}+{sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x}+{sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x}+{sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x}+{sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x}+{sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x}+{sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x}+{sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x}+{sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x}+{sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x}+{sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x}+{sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x}+{sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x}+{sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x}+{sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x}+{sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x}+{sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x}+{sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x}+{sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x}+{sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x}+{sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x}+{sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x}+{sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x}+{sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x}+{sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x}+{sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x}+{sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x}+{sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x}+{sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x}+{sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x}+{sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x}+{sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x}+{sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x}+{sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x}+{sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x}+{sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x}+{sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x}+{sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x}+{sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x}+{sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x}+{sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x}+{sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x}+{sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x}+{sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x}+{sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x}+{sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x}+{sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x}+{sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x}+{sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x}+{sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x}+{sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x}+{sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x}+{sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x}+{sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x}+{sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x}+{sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x}+{sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x}+{sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x}+{sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x}+{sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x}+{sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x}+{sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x}+{sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x}+{sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x}+{sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x}+{sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x}+{sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x}+{sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x}+{sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x}+{sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x}+{sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x}+{sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x}+{sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x}+{sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x}+{sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x}+{sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x}+{sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x}+{sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x}+{sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x}+{sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x}+{sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x}+{sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x}+{sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x}+{sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x}+{sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x}+{sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x}+{sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x}+{sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x}+{sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x}+{sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x}+{sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x}+{sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x}+{sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x}+{sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x}+{sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x}+{sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x}+{sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x}+{B0x[15],B0x[15],B0x[15],B0x[15],B0x[15],B0x[15],B0x[15],B0x};

			if(sumout[22]==0)
				if(sumout[21:13]!=9'b0)
					N1x<=8'd127;
				else
					if(sumout[5]==1 && sumout[4:0]!=5'd0)
						N1x<=sumout[13:6]+8'd1;
					else
						N1x<=sumout[13:6];
			else
				N1x<=8'd0;
			end
		end
endmodule
