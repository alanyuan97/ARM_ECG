module top(EN, clk, reset, out, sel, sel_out);
	input EN, clk, reset;
	output reg [7:0] out;
	input [5:0] sel;
	input [2:0] sel_out;

	wire [1496:0] l1;
	wire [7:0] l2_0, l2_1, l2_2, l2_3, l2_4;
	//wire [7:0] l3_0, l3_1, l3_2, l3_3, l3_4, l3_5, l3_6, l3_7, l3_8, l3_9;
	//wire [7:0] l4_0, l4_1, l4_2, l4_3, l4_4, l4_5, l4_6, l4_7, l4_8, l4_9, l4_10, l4_11, l4_12, l4_13, l4_14;
	//wire [7:0] l5_0, l5_1, l5_2, l5_3, l5_4, l5_5, l5_6, l5_7, l5_8, l5_9, l5_10, l5_11, l5_12, l5_13, l5_14, l5_15, l5_16, l5_17, l5_18, l5_19, l5_20, l5_21, l5_22, l5_23, l5_24, l5_25, l5_26, l5_27, l5_28, l5_29;
	//wire [7:0] l6_0, l6_1, l6_2, l6_3, l6_4, l6_5, l6_6, l6_7, l6_8, l6_9, l6_10, l6_11, l6_12, l6_13, l6_14;
	//wire [7:0] l7_0, l7_1, l7_2, l7_3, l7_4, l7_5, l7_6, l7_7, l7_8, l7_9;


	ROM rom_in(.address(sel),.clock(clk),.q(l1));
	layer_1 layer1(reset, clk, l2_0, l2_1, l2_2, l2_3, l2_4, l1[1495:1488], l1[1487:1480], l1[1479:1472], l1[1471:1464], l1[1463:1456], l1[1455:1448], l1[1447:1440], l1[1439:1432], l1[1431:1424], l1[1423:1416], l1[1415:1408], l1[1407:1400], l1[1399:1392], l1[1391:1384], l1[1383:1376], l1[1375:1368], l1[1367:1360], l1[1359:1352], l1[1351:1344], l1[1343:1336], l1[1335:1328], l1[1327:1320], l1[1319:1312], l1[1311:1304], l1[1303:1296], l1[1295:1288], l1[1287:1280], l1[1279:1272], l1[1271:1264], l1[1263:1256], l1[1255:1248], l1[1247:1240], l1[1239:1232], l1[1231:1224], l1[1223:1216], l1[1215:1208], l1[1207:1200], l1[1199:1192], l1[1191:1184], l1[1183:1176], l1[1175:1168], l1[1167:1160], l1[1159:1152], l1[1151:1144], l1[1143:1136], l1[1135:1128], l1[1127:1120], l1[1119:1112], l1[1111:1104], l1[1103:1096], l1[1095:1088], l1[1087:1080], l1[1079:1072], l1[1071:1064], l1[1063:1056], l1[1055:1048], l1[1047:1040], l1[1039:1032], l1[1031:1024], l1[1023:1016], l1[1015:1008], l1[1007:1000], l1[999:992], l1[991:984], l1[983:976], l1[975:968], l1[967:960], l1[959:952], l1[951:944], l1[943:936], l1[935:928], l1[927:920], l1[919:912], l1[911:904], l1[903:896], l1[895:888], l1[887:880], l1[879:872], l1[871:864], l1[863:856], l1[855:848], l1[847:840], l1[839:832], l1[831:824], l1[823:816], l1[815:808], l1[807:800], l1[799:792], l1[791:784], l1[783:776], l1[775:768], l1[767:760], l1[759:752], l1[751:744], l1[743:736], l1[735:728], l1[727:720], l1[719:712], l1[711:704], l1[703:696], l1[695:688], l1[687:680], l1[679:672], l1[671:664], l1[663:656], l1[655:648], l1[647:640], l1[639:632], l1[631:624], l1[623:616], l1[615:608], l1[607:600], l1[599:592], l1[591:584], l1[583:576], l1[575:568], l1[567:560], l1[559:552], l1[551:544], l1[543:536], l1[535:528], l1[527:520], l1[519:512], l1[511:504], l1[503:496], l1[495:488], l1[487:480], l1[479:472], l1[471:464], l1[463:456], l1[455:448], l1[447:440], l1[439:432], l1[431:424], l1[423:416], l1[415:408], l1[407:400], l1[399:392], l1[391:384], l1[383:376], l1[375:368], l1[367:360], l1[359:352], l1[351:344], l1[343:336], l1[335:328], l1[327:320], l1[319:312], l1[311:304], l1[303:296], l1[295:288], l1[287:280], l1[279:272], l1[271:264], l1[263:256], l1[255:248], l1[247:240], l1[239:232], l1[231:224], l1[223:216], l1[215:208], l1[207:200], l1[199:192], l1[191:184], l1[183:176], l1[175:168], l1[167:160], l1[159:152], l1[151:144], l1[143:136], l1[135:128], l1[127:120], l1[119:112], l1[111:104], l1[103:96], l1[95:88], l1[87:80], l1[79:72], l1[71:64], l1[63:56], l1[55:48], l1[47:40], l1[39:32], l1[31:24], l1[23:16], l1[15:8], l1[7:0]);
	
	always @(*) begin
		case(sel_out)
			3'b000: out<=l2_0;
			3'b001: out<=l2_1;
			3'b010: out<=l2_2;
			3'b011: out<=l2_3;
			3'b100: out<=l2_4;
			default:out<=l2_0;
		endcase
	end
	//layer_2 layer2(reset, clk, l3_0, l3_1, l3_2, l3_3, l3_4, l3_5, l3_6, l3_7, l3_8, l3_9, l2_0, l2_1, l2_2, l2_3, l2_4);
	//layer_3 layer3(reset, clk, l4_0, l4_1, l4_2, l4_3, l4_4, l4_5, l4_6, l4_7, l4_8, l4_9, l4_10, l4_11, l4_12, l4_13, l4_14, l3_0, l3_1, l3_2, l3_3, l3_4, l3_5, l3_6, l3_7, l3_8, l3_9);
	//layer_4 layer4(reset, clk, l5_0, l5_1, l5_2, l5_3, l5_4, l5_5, l5_6, l5_7, l5_8, l5_9, l5_10, l5_11, l5_12, l5_13, l5_14, l5_15, l5_16, l5_17, l5_18, l5_19, l5_20, l5_21, l5_22, l5_23, l5_24, l5_25, l5_26, l5_27, l5_28, l5_29, l4_0, l4_1, l4_2, l4_3, l4_4, l4_5, l4_6, l4_7, l4_8, l4_9, l4_10, l4_11, l4_12, l4_13, l4_14);
	//layer_5 layer5(reset, clk, l6_0, l6_1, l6_2, l6_3, l6_4, l6_5, l6_6, l6_7, l6_8, l6_9, l6_10, l6_11, l6_12, l6_13, l6_14, l5_0, l5_1, l5_2, l5_3, l5_4, l5_5, l5_6, l5_7, l5_8, l5_9, l5_10, l5_11, l5_12, l5_13, l5_14, l5_15, l5_16, l5_17, l5_18, l5_19, l5_20, l5_21, l5_22, l5_23, l5_24, l5_25, l5_26, l5_27, l5_28, l5_29);
	//layer_6 layer6(reset, clk, l7_0, l7_1, l7_2, l7_3, l7_4, l7_5, l7_6, l7_7, l7_8, l7_9, l6_0, l6_1, l6_2, l6_3, l6_4, l6_5, l6_6, l6_7, l6_8, l6_9, l6_10, l6_11, l6_12, l6_13, l6_14);
	//layer_7 layer7(reset, clk, out0, l7_0, l7_1, l7_2, l7_3, l7_4, l7_5, l7_6, l7_7, l7_8, l7_9);
endmodule
