module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 525;
	I1x = 6230;
	I2x = -7406;
	I3x = 1709;
	I4x = 4118;
	I5x = -1828;
	I6x = -2715;
	I7x = 4181;
	I8x = 3276;
	I9x = 1716;
	I10x = -4718;
	I11x = -2391;
	I12x = -1101;
	I13x = -6598;
	I14x = -5481;
	I15x = -849;
	I16x = -413;
	I17x = -3615;
	I18x = -1973;
	I19x = -5139;
	I20x = -1219;
	I21x = -55;
	I22x = 3868;
	I23x = -420;
	I24x = 340;
	I25x = 4094;
	I26x = 0;
	I27x = -6325;
	I28x = 3179;
	I29x = 1675;
	I30x = -7841;
	I31x = -3365;
	I32x = -6011;
	I33x = -65;
	I34x = -174;
	I35x = 5944;
	I36x = -3040;
	I37x = 1864;
	I38x = 2245;
	I39x = 5947;
	I40x = -1372;
	I41x = 1656;
	I42x = -8173;
	I43x = 2444;
	I44x = 1941;
	I45x = -3086;
	I46x = -3378;
	I47x = -5174;
	I48x = 1274;
	I49x = 6264;
	I50x = 2899;
	I51x = 6984;
	I52x = -6934;
	I53x = 7382;
	I54x = 3514;
	I55x = -3178;
	I56x = 3808;
	I57x = -6272;
	I58x = 3346;
	I59x = -391;
	I60x = -2118;
	I61x = 7448;
	I62x = -5172;
	I63x = 2641;
	I64x = 4005;
	I65x = -7137;
	I66x = 4763;
	I67x = 8003;
	I68x = -2154;
	I69x = -2321;
	I70x = -1320;
	I71x = -7644;
	I72x = -5732;
	I73x = 5132;
	I74x = -5708;
	I75x = -5426;
	I76x = -7545;
	I77x = 2519;
	I78x = 4822;
	I79x = -2953;
	I80x = -4365;
	I81x = 5795;
	I82x = -2401;
	I83x = -5538;
	I84x = 5235;
	I85x = 2486;
	I86x = 4414;
	I87x = -5799;
	I88x = -4557;
	I89x = 5681;
	I90x = 2657;
	I91x = -7878;
	I92x = 4400;
	I93x = 1045;
	I94x = -6875;
	I95x = 3182;
	I96x = -5985;
	I97x = -6264;
	I98x = -6310;
	I99x = 5513;
	I100x = 2912;
	I101x = 3434;
	I102x = -4579;
	I103x = -1649;
	I104x = -2787;
	I105x = -5712;
	I106x = -5566;
	I107x = -4296;
	I108x = -7498;
	I109x = -7041;
	I110x = -1340;
	I111x = -2619;
	I112x = 4952;
	I113x = -586;
	I114x = 6574;
	I115x = 3208;
	I116x = -2490;
	I117x = -6250;
	I118x = 1456;
	I119x = -452;
	I120x = -7380;
	I121x = 1780;
	I122x = -6532;
	I123x = 1053;
	I124x = 4599;
	I125x = -4269;
	I126x = -7649;
	I127x = 2530;
	I128x = 2420;
	I129x = 2392;
	I130x = -4717;
	I131x = -2522;
	I132x = 7682;
	I133x = 3454;
	I134x = 7959;
	I135x = 3263;
	I136x = -531;
	I137x = 7060;
	I138x = 5883;
	I139x = 3929;
	I140x = -5738;
	I141x = 7528;
	I142x = -1157;
	I143x = 1704;
	I144x = 4971;
	I145x = -6651;
	I146x = 5699;
	I147x = 2805;
	I148x = 7482;
	I149x = -4360;
	I150x = -4658;
	I151x = 4500;
	I152x = -679;
	I153x = 5769;
	I154x = -91;
	I155x = -4981;
	I156x = -2230;
	I157x = -4640;
	I158x = 1143;
	I159x = -3858;
	I160x = 127;
	I161x = -2855;
	I162x = -6999;
	I163x = 3912;
	I164x = 5187;
	I165x = 3367;
	I166x = -63;
	I167x = -1249;
	I168x = -6254;
	I169x = -2051;
	I170x = -5452;
	I171x = 8062;
	I172x = 1450;
	I173x = 2021;
	I174x = 1332;
	I175x = -5696;
	I176x = -8165;
	I177x = -233;
	I178x = 5608;
	I179x = -5271;
	I180x = 7493;
	I181x = 5824;
	I182x = -257;
	I183x = -2987;
	I184x = -5747;
	I185x = 5599;
	I186x = 2591;
	end
endmodule
[2.7983595  0.         0.         0.25730097 0.        ] 

 [22924, 0, 0, 2107, 0] 

 ['0101100110001100', '0000000000000000', '0000000000000000', '0000100000111011', '0000000000000000']
