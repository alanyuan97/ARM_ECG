module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 7355;
	I1x = 639;
	I2x = -1996;
	I3x = -1755;
	I4x = 3671;
	I5x = 1319;
	I6x = -7014;
	I7x = -6603;
	I8x = -2466;
	I9x = 3200;
	I10x = 4150;
	I11x = -7284;
	I12x = 7404;
	I13x = 5695;
	I14x = 5320;
	I15x = -4349;
	I16x = -5913;
	I17x = 8183;
	I18x = 3792;
	I19x = -2540;
	I20x = -3399;
	I21x = -734;
	I22x = -3888;
	I23x = -3611;
	I24x = -4078;
	I25x = 4789;
	I26x = 3906;
	I27x = 488;
	I28x = -4698;
	I29x = 7634;
	I30x = -4710;
	I31x = -433;
	I32x = 3085;
	I33x = 3506;
	I34x = 5763;
	I35x = -5825;
	I36x = 7037;
	I37x = -7702;
	I38x = 4129;
	I39x = 3923;
	I40x = -5042;
	I41x = -3263;
	I42x = -379;
	I43x = -902;
	I44x = -7069;
	I45x = 3725;
	I46x = 615;
	I47x = 3542;
	I48x = 5597;
	I49x = -6592;
	I50x = 5717;
	I51x = 529;
	I52x = -2161;
	I53x = 7341;
	I54x = 3484;
	I55x = -3414;
	I56x = -1576;
	I57x = -1009;
	I58x = -6029;
	I59x = -6746;
	I60x = -4037;
	I61x = 2030;
	I62x = 5750;
	I63x = -6271;
	I64x = 3671;
	I65x = -2460;
	I66x = -5515;
	I67x = 6563;
	I68x = 3322;
	I69x = 2509;
	I70x = -7347;
	I71x = 3684;
	I72x = 7434;
	I73x = -6257;
	I74x = 7305;
	I75x = 4540;
	I76x = 1104;
	I77x = -1626;
	I78x = 1019;
	I79x = -5628;
	I80x = -3009;
	I81x = 6200;
	I82x = -1588;
	I83x = -1358;
	I84x = -1309;
	I85x = -4005;
	I86x = -5124;
	I87x = 6411;
	I88x = -4106;
	I89x = -7938;
	I90x = 2249;
	I91x = -6466;
	I92x = 2965;
	I93x = 8118;
	I94x = -4506;
	I95x = 6781;
	I96x = 1004;
	I97x = 1567;
	I98x = 5916;
	I99x = 3688;
	I100x = -1931;
	I101x = -4966;
	I102x = 7533;
	I103x = 3213;
	I104x = -3110;
	I105x = -1348;
	I106x = -6271;
	I107x = -6356;
	I108x = 885;
	I109x = 2483;
	I110x = 6034;
	I111x = -7712;
	I112x = -7245;
	I113x = 1400;
	I114x = 803;
	I115x = 1715;
	I116x = 2152;
	I117x = 2882;
	I118x = 3512;
	I119x = -4423;
	I120x = 4308;
	I121x = -253;
	I122x = -4961;
	I123x = 7526;
	I124x = 6016;
	I125x = 3589;
	I126x = 3011;
	I127x = -7630;
	I128x = 3000;
	I129x = -4055;
	I130x = 502;
	I131x = -1130;
	I132x = -498;
	I133x = -7694;
	I134x = 8147;
	I135x = -5579;
	I136x = -5543;
	I137x = -5614;
	I138x = -1684;
	I139x = -6188;
	I140x = -1016;
	I141x = -564;
	I142x = 4514;
	I143x = -2993;
	I144x = 3418;
	I145x = -7750;
	I146x = -1392;
	I147x = 6038;
	I148x = -1324;
	I149x = -6288;
	I150x = 4085;
	I151x = -5086;
	I152x = -6635;
	I153x = -5846;
	I154x = -3843;
	I155x = -7330;
	I156x = -8052;
	I157x = -4212;
	I158x = 1979;
	I159x = 6266;
	I160x = -398;
	I161x = -4595;
	I162x = 8151;
	I163x = 3856;
	I164x = 2096;
	I165x = 5942;
	I166x = -5130;
	I167x = 204;
	I168x = -5257;
	I169x = -2112;
	I170x = 5437;
	I171x = 4046;
	I172x = 4012;
	I173x = -6742;
	I174x = -2032;
	I175x = 4091;
	I176x = -1951;
	I177x = 5239;
	I178x = 7521;
	I179x = 5870;
	I180x = -2265;
	I181x = 971;
	I182x = -7773;
	I183x = 4398;
	I184x = -2027;
	I185x = 6447;
	I186x = -5750;
	end
endmodule
[1.05815576 0.35814832 2.61052972 0.         0.45510654] 

 [8668, 2933, 21385, 0, 3728] 

 ['0010000111011100', '0000101101110101', '0101001110001001', '0000000000000000', '0000111010010000']
