module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 5189;
	I1x = -1406;
	I2x = 1599;
	I3x = -5759;
	I4x = 7304;
	I5x = 4076;
	I6x = 4523;
	I7x = -3870;
	I8x = 2081;
	I9x = 2872;
	I10x = 1359;
	I11x = -7436;
	I12x = 3280;
	I13x = -1931;
	I14x = 8154;
	I15x = 2698;
	I16x = -3548;
	I17x = 5349;
	I18x = -3497;
	I19x = 3059;
	I20x = -6584;
	I21x = 5006;
	I22x = -4281;
	I23x = -8057;
	I24x = -3874;
	I25x = 3115;
	I26x = 472;
	I27x = 3125;
	I28x = -2775;
	I29x = -7535;
	I30x = 7923;
	I31x = -7211;
	I32x = -4266;
	I33x = -5186;
	I34x = -2852;
	I35x = -6026;
	I36x = 7658;
	I37x = 1392;
	I38x = 6743;
	I39x = 3854;
	I40x = 2162;
	I41x = -815;
	I42x = -6752;
	I43x = -6213;
	I44x = -4;
	I45x = -7057;
	I46x = -3634;
	I47x = -7625;
	I48x = -3154;
	I49x = 3562;
	I50x = -7127;
	I51x = 7536;
	I52x = 608;
	I53x = 7194;
	I54x = -6796;
	I55x = 399;
	I56x = -6234;
	I57x = 7129;
	I58x = -6250;
	I59x = -1042;
	I60x = -4971;
	I61x = 149;
	I62x = -5954;
	I63x = -678;
	I64x = 2648;
	I65x = -5014;
	I66x = -3154;
	I67x = -5478;
	I68x = 3584;
	I69x = 1862;
	I70x = 7767;
	I71x = -4869;
	I72x = -2034;
	I73x = 7308;
	I74x = 2079;
	I75x = -6883;
	I76x = -7931;
	I77x = -1684;
	I78x = 6378;
	I79x = -1067;
	I80x = 2246;
	I81x = 333;
	I82x = 6937;
	I83x = -2037;
	I84x = 2438;
	I85x = -6328;
	I86x = 1868;
	I87x = 7815;
	I88x = -3548;
	I89x = 5418;
	I90x = 6669;
	I91x = 6919;
	I92x = -6471;
	I93x = 6687;
	I94x = 3936;
	I95x = -5157;
	I96x = 6406;
	I97x = -2801;
	I98x = -1156;
	I99x = 6635;
	I100x = 8031;
	I101x = 5947;
	I102x = -2107;
	I103x = -465;
	I104x = 5720;
	I105x = 6835;
	I106x = -912;
	I107x = 4172;
	I108x = 7228;
	I109x = -3086;
	I110x = 566;
	I111x = 3899;
	I112x = -5420;
	I113x = -124;
	I114x = -1439;
	I115x = 4081;
	I116x = 5009;
	I117x = -4217;
	I118x = 6498;
	I119x = -3976;
	I120x = -3019;
	I121x = -53;
	I122x = 6558;
	I123x = 600;
	I124x = 2332;
	I125x = 1799;
	I126x = 2778;
	I127x = -2430;
	I128x = 6270;
	I129x = -4730;
	I130x = -3999;
	I131x = 7220;
	I132x = 843;
	I133x = 1648;
	I134x = 7411;
	I135x = 1019;
	I136x = -7533;
	I137x = -2802;
	I138x = -712;
	I139x = -4707;
	I140x = -5274;
	I141x = 7186;
	I142x = -8001;
	I143x = 1010;
	I144x = -1659;
	I145x = -3331;
	I146x = -7212;
	I147x = 1687;
	I148x = -2267;
	I149x = -6607;
	I150x = 3760;
	I151x = 5130;
	I152x = 4175;
	I153x = -1071;
	I154x = 7259;
	I155x = 2283;
	I156x = 1750;
	I157x = -2313;
	I158x = 1181;
	I159x = 1987;
	I160x = -3760;
	I161x = 8027;
	I162x = 6686;
	I163x = 2306;
	I164x = -4022;
	I165x = 4122;
	I166x = 1071;
	I167x = 754;
	I168x = 3206;
	I169x = 2102;
	I170x = 8182;
	I171x = -4803;
	I172x = -2964;
	I173x = 1386;
	I174x = -4165;
	I175x = -4098;
	I176x = -60;
	I177x = -4455;
	I178x = -1087;
	I179x = -4894;
	I180x = 6443;
	I181x = 3226;
	I182x = -7920;
	I183x = 170;
	I184x = -4987;
	I185x = -749;
	I186x = -6226;
	end
endmodule
[0.02602729 0.         0.         0.         0.        ] 

 [213, 0, 0, 0, 0] 

 ['0000000011010101', '0000000000000000', '0000000000000000', '0000000000000000', '0000000000000000']
