module top(EN, clk, reset, out0);
	input EN, clk, reset;
	output [7:0] out0;

	wire [7:0] l1_0, l1_1, l1_2, l1_3, l1_4, l1_5, l1_6, l1_7, l1_8, l1_9, l1_10, l1_11, l1_12, l1_13, l1_14, l1_15, l1_16, l1_17, l1_18, l1_19, l1_20, l1_21, l1_22, l1_23, l1_24, l1_25, l1_26, l1_27, l1_28, l1_29, l1_30, l1_31, l1_32, l1_33, l1_34, l1_35, l1_36, l1_37, l1_38, l1_39, l1_40, l1_41, l1_42, l1_43, l1_44, l1_45, l1_46, l1_47, l1_48, l1_49, l1_50, l1_51, l1_52, l1_53, l1_54, l1_55, l1_56, l1_57, l1_58, l1_59, l1_60, l1_61, l1_62, l1_63, l1_64, l1_65, l1_66, l1_67, l1_68, l1_69, l1_70, l1_71, l1_72, l1_73, l1_74, l1_75, l1_76, l1_77, l1_78, l1_79, l1_80, l1_81, l1_82, l1_83, l1_84, l1_85, l1_86, l1_87, l1_88, l1_89, l1_90, l1_91, l1_92, l1_93, l1_94, l1_95, l1_96, l1_97, l1_98, l1_99, l1_100, l1_101, l1_102, l1_103, l1_104, l1_105, l1_106, l1_107, l1_108, l1_109, l1_110, l1_111, l1_112, l1_113, l1_114, l1_115, l1_116, l1_117, l1_118, l1_119, l1_120, l1_121, l1_122, l1_123, l1_124, l1_125, l1_126, l1_127, l1_128, l1_129, l1_130, l1_131, l1_132, l1_133, l1_134, l1_135, l1_136, l1_137, l1_138, l1_139, l1_140, l1_141, l1_142, l1_143, l1_144, l1_145, l1_146, l1_147, l1_148, l1_149, l1_150, l1_151, l1_152, l1_153, l1_154, l1_155, l1_156, l1_157, l1_158, l1_159, l1_160, l1_161, l1_162, l1_163, l1_164, l1_165, l1_166, l1_167, l1_168, l1_169, l1_170, l1_171, l1_172, l1_173, l1_174, l1_175, l1_176, l1_177, l1_178, l1_179, l1_180, l1_181, l1_182, l1_183, l1_184, l1_185, l1_186;
	wire [7:0] l2_0, l2_1, l2_2, l2_3, l2_4;
	wire [7:0] l3_0, l3_1, l3_2, l3_3, l3_4, l3_5, l3_6, l3_7, l3_8, l3_9;
	wire [7:0] l4_0, l4_1, l4_2, l4_3, l4_4, l4_5, l4_6, l4_7, l4_8, l4_9, l4_10, l4_11, l4_12, l4_13, l4_14;
	wire [7:0] l5_0, l5_1, l5_2, l5_3, l5_4, l5_5, l5_6, l5_7, l5_8, l5_9, l5_10, l5_11, l5_12, l5_13, l5_14, l5_15, l5_16, l5_17, l5_18, l5_19, l5_20, l5_21, l5_22, l5_23, l5_24, l5_25, l5_26, l5_27, l5_28, l5_29;
	wire [7:0] l6_0, l6_1, l6_2, l6_3, l6_4, l6_5, l6_6, l6_7, l6_8, l6_9, l6_10, l6_11, l6_12, l6_13, l6_14;
	wire [7:0] l7_0, l7_1, l7_2, l7_3, l7_4, l7_5, l7_6, l7_7, l7_8, l7_9;


	rom_input rom_in(EN, clk, l1_0, l1_1, l1_2, l1_3, l1_4, l1_5, l1_6, l1_7, l1_8, l1_9, l1_10, l1_11, l1_12, l1_13, l1_14, l1_15, l1_16, l1_17, l1_18, l1_19, l1_20, l1_21, l1_22, l1_23, l1_24, l1_25, l1_26, l1_27, l1_28, l1_29, l1_30, l1_31, l1_32, l1_33, l1_34, l1_35, l1_36, l1_37, l1_38, l1_39, l1_40, l1_41, l1_42, l1_43, l1_44, l1_45, l1_46, l1_47, l1_48, l1_49, l1_50, l1_51, l1_52, l1_53, l1_54, l1_55, l1_56, l1_57, l1_58, l1_59, l1_60, l1_61, l1_62, l1_63, l1_64, l1_65, l1_66, l1_67, l1_68, l1_69, l1_70, l1_71, l1_72, l1_73, l1_74, l1_75, l1_76, l1_77, l1_78, l1_79, l1_80, l1_81, l1_82, l1_83, l1_84, l1_85, l1_86, l1_87, l1_88, l1_89, l1_90, l1_91, l1_92, l1_93, l1_94, l1_95, l1_96, l1_97, l1_98, l1_99, l1_100, l1_101, l1_102, l1_103, l1_104, l1_105, l1_106, l1_107, l1_108, l1_109, l1_110, l1_111, l1_112, l1_113, l1_114, l1_115, l1_116, l1_117, l1_118, l1_119, l1_120, l1_121, l1_122, l1_123, l1_124, l1_125, l1_126, l1_127, l1_128, l1_129, l1_130, l1_131, l1_132, l1_133, l1_134, l1_135, l1_136, l1_137, l1_138, l1_139, l1_140, l1_141, l1_142, l1_143, l1_144, l1_145, l1_146, l1_147, l1_148, l1_149, l1_150, l1_151, l1_152, l1_153, l1_154, l1_155, l1_156, l1_157, l1_158, l1_159, l1_160, l1_161, l1_162, l1_163, l1_164, l1_165, l1_166, l1_167, l1_168, l1_169, l1_170, l1_171, l1_172, l1_173, l1_174, l1_175, l1_176, l1_177, l1_178, l1_179, l1_180, l1_181, l1_182, l1_183, l1_184, l1_185, l1_186);
	layer_1 layer1(reset, clk, l2_0, l2_1, l2_2, l2_3, l2_4, l1_0, l1_1, l1_2, l1_3, l1_4, l1_5, l1_6, l1_7, l1_8, l1_9, l1_10, l1_11, l1_12, l1_13, l1_14, l1_15, l1_16, l1_17, l1_18, l1_19, l1_20, l1_21, l1_22, l1_23, l1_24, l1_25, l1_26, l1_27, l1_28, l1_29, l1_30, l1_31, l1_32, l1_33, l1_34, l1_35, l1_36, l1_37, l1_38, l1_39, l1_40, l1_41, l1_42, l1_43, l1_44, l1_45, l1_46, l1_47, l1_48, l1_49, l1_50, l1_51, l1_52, l1_53, l1_54, l1_55, l1_56, l1_57, l1_58, l1_59, l1_60, l1_61, l1_62, l1_63, l1_64, l1_65, l1_66, l1_67, l1_68, l1_69, l1_70, l1_71, l1_72, l1_73, l1_74, l1_75, l1_76, l1_77, l1_78, l1_79, l1_80, l1_81, l1_82, l1_83, l1_84, l1_85, l1_86, l1_87, l1_88, l1_89, l1_90, l1_91, l1_92, l1_93, l1_94, l1_95, l1_96, l1_97, l1_98, l1_99, l1_100, l1_101, l1_102, l1_103, l1_104, l1_105, l1_106, l1_107, l1_108, l1_109, l1_110, l1_111, l1_112, l1_113, l1_114, l1_115, l1_116, l1_117, l1_118, l1_119, l1_120, l1_121, l1_122, l1_123, l1_124, l1_125, l1_126, l1_127, l1_128, l1_129, l1_130, l1_131, l1_132, l1_133, l1_134, l1_135, l1_136, l1_137, l1_138, l1_139, l1_140, l1_141, l1_142, l1_143, l1_144, l1_145, l1_146, l1_147, l1_148, l1_149, l1_150, l1_151, l1_152, l1_153, l1_154, l1_155, l1_156, l1_157, l1_158, l1_159, l1_160, l1_161, l1_162, l1_163, l1_164, l1_165, l1_166, l1_167, l1_168, l1_169, l1_170, l1_171, l1_172, l1_173, l1_174, l1_175, l1_176, l1_177, l1_178, l1_179, l1_180, l1_181, l1_182, l1_183, l1_184, l1_185, l1_186);
	layer_2 layer2(reset, clk, l3_0, l3_1, l3_2, l3_3, l3_4, l3_5, l3_6, l3_7, l3_8, l3_9, l2_0, l2_1, l2_2, l2_3, l2_4);
	layer_3 layer3(reset, clk, l4_0, l4_1, l4_2, l4_3, l4_4, l4_5, l4_6, l4_7, l4_8, l4_9, l4_10, l4_11, l4_12, l4_13, l4_14, l3_0, l3_1, l3_2, l3_3, l3_4, l3_5, l3_6, l3_7, l3_8, l3_9);
	layer_4 layer4(reset, clk, l5_0, l5_1, l5_2, l5_3, l5_4, l5_5, l5_6, l5_7, l5_8, l5_9, l5_10, l5_11, l5_12, l5_13, l5_14, l5_15, l5_16, l5_17, l5_18, l5_19, l5_20, l5_21, l5_22, l5_23, l5_24, l5_25, l5_26, l5_27, l5_28, l5_29, l4_0, l4_1, l4_2, l4_3, l4_4, l4_5, l4_6, l4_7, l4_8, l4_9, l4_10, l4_11, l4_12, l4_13, l4_14);
	layer_5 layer5(reset, clk, l6_0, l6_1, l6_2, l6_3, l6_4, l6_5, l6_6, l6_7, l6_8, l6_9, l6_10, l6_11, l6_12, l6_13, l6_14, l5_0, l5_1, l5_2, l5_3, l5_4, l5_5, l5_6, l5_7, l5_8, l5_9, l5_10, l5_11, l5_12, l5_13, l5_14, l5_15, l5_16, l5_17, l5_18, l5_19, l5_20, l5_21, l5_22, l5_23, l5_24, l5_25, l5_26, l5_27, l5_28, l5_29);
	layer_6 layer6(reset, clk, l7_0, l7_1, l7_2, l7_3, l7_4, l7_5, l7_6, l7_7, l7_8, l7_9, l6_0, l6_1, l6_2, l6_3, l6_4, l6_5, l6_6, l6_7, l6_8, l6_9, l6_10, l6_11, l6_12, l6_13, l6_14);
	layer_7 layer7(reset, clk, out0, l7_0, l7_1, l7_2, l7_3, l7_4, l7_5, l7_6, l7_7, l7_8, l7_9);
endmodule
