module node1_5(N1A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,A16,A17,A18,A19,A20,A21,A22,A23,A24,A25,A26,A27,A28,A29,A30,A31,A32,A33,A34,A35,A36,A37,A38,A39,A40,A41,A42,A43,A44,A45,A46,A47,A48,A49,A50,A51,A52,A53,A54,A55,A56,A57,A58,A59,A60,A61,A62,A63,A64,A65,A66,A67,A68,A69,A70,A71,A72,A73,A74,A75,A76,A77,A78,A79,A80,A81,A82,A83,A84,A85,A86,A87,A88,A89,A90,A91,A92,A93,A94,A95,A96,A97,A98,A99,A100,A101,A102,A103,A104,A105,A106,A107,A108,A109,A110,A111,A112,A113,A114,A115,A116,A117,A118,A119,A120,A121,A122,A123,A124,A125,A126,A127,A128,A129,A130,A131,A132,A133,A134,A135,A136,A137,A138,A139,A140,A141,A142,A143,A144,A145,A146,A147,A148,A149,A150,A151,A152,A153,A154,A155,A156,A157,A158,A159,A160,A161,A162,A163,A164,A165,A166,A167,A168,A169,A170,A171,A172,A173,A174,A175,A176,A177,A178,A179,A180,A181,A182,A183,A184,A185,A186);
	input [31:0] A0;
	input [31:0] A1;
	input [31:0] A2;
	input [31:0] A3;
	input [31:0] A4;
	input [31:0] A5;
	input [31:0] A6;
	input [31:0] A7;
	input [31:0] A8;
	input [31:0] A9;
	input [31:0] A10;
	input [31:0] A11;
	input [31:0] A12;
	input [31:0] A13;
	input [31:0] A14;
	input [31:0] A15;
	input [31:0] A16;
	input [31:0] A17;
	input [31:0] A18;
	input [31:0] A19;
	input [31:0] A20;
	input [31:0] A21;
	input [31:0] A22;
	input [31:0] A23;
	input [31:0] A24;
	input [31:0] A25;
	input [31:0] A26;
	input [31:0] A27;
	input [31:0] A28;
	input [31:0] A29;
	input [31:0] A30;
	input [31:0] A31;
	input [31:0] A32;
	input [31:0] A33;
	input [31:0] A34;
	input [31:0] A35;
	input [31:0] A36;
	input [31:0] A37;
	input [31:0] A38;
	input [31:0] A39;
	input [31:0] A40;
	input [31:0] A41;
	input [31:0] A42;
	input [31:0] A43;
	input [31:0] A44;
	input [31:0] A45;
	input [31:0] A46;
	input [31:0] A47;
	input [31:0] A48;
	input [31:0] A49;
	input [31:0] A50;
	input [31:0] A51;
	input [31:0] A52;
	input [31:0] A53;
	input [31:0] A54;
	input [31:0] A55;
	input [31:0] A56;
	input [31:0] A57;
	input [31:0] A58;
	input [31:0] A59;
	input [31:0] A60;
	input [31:0] A61;
	input [31:0] A62;
	input [31:0] A63;
	input [31:0] A64;
	input [31:0] A65;
	input [31:0] A66;
	input [31:0] A67;
	input [31:0] A68;
	input [31:0] A69;
	input [31:0] A70;
	input [31:0] A71;
	input [31:0] A72;
	input [31:0] A73;
	input [31:0] A74;
	input [31:0] A75;
	input [31:0] A76;
	input [31:0] A77;
	input [31:0] A78;
	input [31:0] A79;
	input [31:0] A80;
	input [31:0] A81;
	input [31:0] A82;
	input [31:0] A83;
	input [31:0] A84;
	input [31:0] A85;
	input [31:0] A86;
	input [31:0] A87;
	input [31:0] A88;
	input [31:0] A89;
	input [31:0] A90;
	input [31:0] A91;
	input [31:0] A92;
	input [31:0] A93;
	input [31:0] A94;
	input [31:0] A95;
	input [31:0] A96;
	input [31:0] A97;
	input [31:0] A98;
	input [31:0] A99;
	input [31:0] A100;
	input [31:0] A101;
	input [31:0] A102;
	input [31:0] A103;
	input [31:0] A104;
	input [31:0] A105;
	input [31:0] A106;
	input [31:0] A107;
	input [31:0] A108;
	input [31:0] A109;
	input [31:0] A110;
	input [31:0] A111;
	input [31:0] A112;
	input [31:0] A113;
	input [31:0] A114;
	input [31:0] A115;
	input [31:0] A116;
	input [31:0] A117;
	input [31:0] A118;
	input [31:0] A119;
	input [31:0] A120;
	input [31:0] A121;
	input [31:0] A122;
	input [31:0] A123;
	input [31:0] A124;
	input [31:0] A125;
	input [31:0] A126;
	input [31:0] A127;
	input [31:0] A128;
	input [31:0] A129;
	input [31:0] A130;
	input [31:0] A131;
	input [31:0] A132;
	input [31:0] A133;
	input [31:0] A134;
	input [31:0] A135;
	input [31:0] A136;
	input [31:0] A137;
	input [31:0] A138;
	input [31:0] A139;
	input [31:0] A140;
	input [31:0] A141;
	input [31:0] A142;
	input [31:0] A143;
	input [31:0] A144;
	input [31:0] A145;
	input [31:0] A146;
	input [31:0] A147;
	input [31:0] A148;
	input [31:0] A149;
	input [31:0] A150;
	input [31:0] A151;
	input [31:0] A152;
	input [31:0] A153;
	input [31:0] A154;
	input [31:0] A155;
	input [31:0] A156;
	input [31:0] A157;
	input [31:0] A158;
	input [31:0] A159;
	input [31:0] A160;
	input [31:0] A161;
	input [31:0] A162;
	input [31:0] A163;
	input [31:0] A164;
	input [31:0] A165;
	input [31:0] A166;
	input [31:0] A167;
	input [31:0] A168;
	input [31:0] A169;
	input [31:0] A170;
	input [31:0] A171;
	input [31:0] A172;
	input [31:0] A173;
	input [31:0] A174;
	input [31:0] A175;
	input [31:0] A176;
	input [31:0] A177;
	input [31:0] A178;
	input [31:0] A179;
	input [31:0] A180;
	input [31:0] A181;
	input [31:0] A182;
	input [31:0] A183;
	input [31:0] A184;
	input [31:0] A185;
	input [31:0] A186;
	output [31:0] N1;

	parameter [31:0] W0=32'b00111101110110010101110110011111;
	parameter [31:0] W1=32'b00111100111110001101011101101110;
	parameter [31:0] W2=32'b10111100111101111010111011001000;
	parameter [31:0] W3=32'b00111110001111110100001010101011;
	parameter [31:0] W4=32'b00111101100001001001110000101010;
	parameter [31:0] W5=32'b00111101110101001111101010111001;
	parameter [31:0] W6=32'b00111101000111011100101100010010;
	parameter [31:0] W7=32'b10111100100010001010001101100100;
	parameter [31:0] W8=32'b10111101011111011101110011010001;
	parameter [31:0] W9=32'b00111101110101111101111100001011;
	parameter [31:0] W10=32'b10111101110111011111000011001010;
	parameter [31:0] W11=32'b00111110010110010100100110100011;
	parameter [31:0] W12=32'b00111110010000001011001010111010;
	parameter [31:0] W13=32'b00111101000000110101010000100111;
	parameter [31:0] W14=32'b00111110010011111101000000100000;
	parameter [31:0] W15=32'b00111110100111100111111110000110;
	parameter [31:0] W16=32'b00111110011100001000000001110011;
	parameter [31:0] W17=32'b00111110101101010010111101001011;
	parameter [31:0] W18=32'b10111011011100100100001011110100;
	parameter [31:0] W19=32'b00111101111001011111111110000000;
	parameter [31:0] W20=32'b10111101010011100000111011000100;
	parameter [31:0] W21=32'b10111101001101011100101100111111;
	parameter [31:0] W22=32'b00111110000101100001010110011101;
	parameter [31:0] W23=32'b10111110010110010000101000001011;
	parameter [31:0] W24=32'b10111101101111101010010010101001;
	parameter [31:0] W25=32'b10111110100100010000000001100010;
	parameter [31:0] W26=32'b10111110100111100110110101010011;
	parameter [31:0] W27=32'b10111110010010110110000111010101;
	parameter [31:0] W28=32'b10111110111000110111110111100001;
	parameter [31:0] W29=32'b10111110111110001101010110010100;
	parameter [31:0] W30=32'b10111110110101011110110001110111;
	parameter [31:0] W31=32'b10111110110110010001101000100011;
	parameter [31:0] W32=32'b10111110101010011110000110101011;
	parameter [31:0] W33=32'b10111110100100010000110011100100;
	parameter [31:0] W34=32'b10111100101000101100001100111000;
	parameter [31:0] W35=32'b00111110000101110100010100100010;
	parameter [31:0] W36=32'b00111110101100100111001010011101;
	parameter [31:0] W37=32'b00111110110111000000111110111011;
	parameter [31:0] W38=32'b00111101111010000011100110101111;
	parameter [31:0] W39=32'b00111101010011111010011100111010;
	parameter [31:0] W40=32'b00111110010110001001011000110100;
	parameter [31:0] W41=32'b00111110000110110001010101110101;
	parameter [31:0] W42=32'b10111110000101010011010111100110;
	parameter [31:0] W43=32'b10111100110110100001110111100100;
	parameter [31:0] W44=32'b10111100111111100110101010101110;
	parameter [31:0] W45=32'b10111101100000110000010010011010;
	parameter [31:0] W46=32'b00111101100010110100111010010111;
	parameter [31:0] W47=32'b00111100100101001000010111010111;
	parameter [31:0] W48=32'b10111011100100010110000010000101;
	parameter [31:0] W49=32'b00111101010110100100101101010100;
	parameter [31:0] W50=32'b00111110011110000110100101010101;
	parameter [31:0] W51=32'b00111110001011000010100001100101;
	parameter [31:0] W52=32'b10111101110101100010101001111000;
	parameter [31:0] W53=32'b10111101110101001100100011100010;
	parameter [31:0] W54=32'b10111101011010101011011000000011;
	parameter [31:0] W55=32'b00111110000101010010001101001100;
	parameter [31:0] W56=32'b00111110001100010011000011100111;
	parameter [31:0] W57=32'b00111110001011101100011111101100;
	parameter [31:0] W58=32'b00111101111100100111011000111011;
	parameter [31:0] W59=32'b00111110100001111010010011010110;
	parameter [31:0] W60=32'b00111110000101000011100000111010;
	parameter [31:0] W61=32'b00111101111001101010010001001001;
	parameter [31:0] W62=32'b00111100100011011010010100110001;
	parameter [31:0] W63=32'b00111110000110111110000101011100;
	parameter [31:0] W64=32'b00111101100001011111101011011100;
	parameter [31:0] W65=32'b00111100100111001000100011001011;
	parameter [31:0] W66=32'b00111110000101110000110110001001;
	parameter [31:0] W67=32'b00111110010000001011111010100001;
	parameter [31:0] W68=32'b10111110000000001010010010001111;
	parameter [31:0] W69=32'b00111101010000100000101011101111;
	parameter [31:0] W70=32'b10111101011110001111101010011010;
	parameter [31:0] W71=32'b10111110100001001110110100100111;
	parameter [31:0] W72=32'b10111110001010010001100001000011;
	parameter [31:0] W73=32'b10111101011111010111101000010110;
	parameter [31:0] W74=32'b10111101000011111110000011110100;
	parameter [31:0] W75=32'b10111100000001000110110100110101;
	parameter [31:0] W76=32'b00111101000100001101111000001000;
	parameter [31:0] W77=32'b00111011100001100110111001010101;
	parameter [31:0] W78=32'b00111011000111110011000100110101;
	parameter [31:0] W79=32'b10111101100101010011010011000100;
	parameter [31:0] W80=32'b00111101001000111001000010101110;
	parameter [31:0] W81=32'b00111101100011010010011100101101;
	parameter [31:0] W82=32'b00111110000001100000000010011010;
	parameter [31:0] W83=32'b10111101100000000100101011000010;
	parameter [31:0] W84=32'b00111101000101101010000000001110;
	parameter [31:0] W85=32'b10111100001110010111101110110010;
	parameter [31:0] W86=32'b00111101111110111101011111111111;
	parameter [31:0] W87=32'b00111100110001101110100010111010;
	parameter [31:0] W88=32'b00111101101001101001111001010100;
	parameter [31:0] W89=32'b00111100100111100101110101001110;
	parameter [31:0] W90=32'b00111101011101000000010000010011;
	parameter [31:0] W91=32'b10111100010000110010100011011110;
	parameter [31:0] W92=32'b00111101110010110001100111010001;
	parameter [31:0] W93=32'b10111100100101110011001001001110;
	parameter [31:0] W94=32'b00111100010001110111000100100010;
	parameter [31:0] W95=32'b00111101100010101111000101011010;
	parameter [31:0] W96=32'b00111101011000010101110011100101;
	parameter [31:0] W97=32'b00111100010011110100011011001011;
	parameter [31:0] W98=32'b10111011001001011010110000100010;
	parameter [31:0] W99=32'b00111100100010010011101110010010;
	parameter [31:0] W100=32'b00111101111011110001110101011000;
	parameter [31:0] W101=32'b10111100101100010010101100011111;
	parameter [31:0] W102=32'b00111101111001000101110110011010;
	parameter [31:0] W103=32'b10111101011101011010110101000101;
	parameter [31:0] W104=32'b00111100100100100011101100010101;
	parameter [31:0] W105=32'b00111101001110011000010100110110;
	parameter [31:0] W106=32'b00111101000110110011011000000000;
	parameter [31:0] W107=32'b00111101001110100111010001001100;
	parameter [31:0] W108=32'b10111110000111111110101110111001;
	parameter [31:0] W109=32'b10111101101000111111110111111101;
	parameter [31:0] W110=32'b00111101010110100001110001010101;
	parameter [31:0] W111=32'b00111100010000000111010011001001;
	parameter [31:0] W112=32'b10111110100100001111010001011100;
	parameter [31:0] W113=32'b10111100011100000110111100011000;
	parameter [31:0] W114=32'b10111101101110111001100001001001;
	parameter [31:0] W115=32'b00111101110001101001000010110111;
	parameter [31:0] W116=32'b10111101010000111101100000001100;
	parameter [31:0] W117=32'b10111101100011000111100000000101;
	parameter [31:0] W118=32'b00111101100111001111100000001101;
	parameter [31:0] W119=32'b10111110100110100100100101010100;
	parameter [31:0] W120=32'b10111110000010101000100110000000;
	parameter [31:0] W121=32'b00111101001100100111001110011100;
	parameter [31:0] W122=32'b00111101001101010001110110000011;
	parameter [31:0] W123=32'b10111101111011011001000110011011;
	parameter [31:0] W124=32'b00111100011010011000010011101111;
	parameter [31:0] W125=32'b10111101110110011011010111010100;
	parameter [31:0] W126=32'b00111100000000111100100000011100;
	parameter [31:0] W127=32'b00111101001101110011110111110000;
	parameter [31:0] W128=32'b10111101000001000111100001001010;
	parameter [31:0] W129=32'b10111110100000111100111101000111;
	parameter [31:0] W130=32'b10111110000011000111011101000111;
	parameter [31:0] W131=32'b10111110101011110100101001101101;
	parameter [31:0] W132=32'b10111110011010011100101011010011;
	parameter [31:0] W133=32'b10111110001000101110010000100011;
	parameter [31:0] W134=32'b10111110100101001011110001101001;
	parameter [31:0] W135=32'b10111110000001111110110010001010;
	parameter [31:0] W136=32'b10111110011000110000001100010000;
	parameter [31:0] W137=32'b10111110001110101010101111101001;
	parameter [31:0] W138=32'b10111110110000111000111001101101;
	parameter [31:0] W139=32'b10111101110000001011110111101100;
	parameter [31:0] W140=32'b10111110001011000100011001101010;
	parameter [31:0] W141=32'b00111101110000100100100001101010;
	parameter [31:0] W142=32'b10111110100001001100101101011100;
	parameter [31:0] W143=32'b00111100101101110110011111011111;
	parameter [31:0] W144=32'b00111101000110001101001100010001;
	parameter [31:0] W145=32'b10111011110111111111011011110000;
	parameter [31:0] W146=32'b10111101100011110001010110010010;
	parameter [31:0] W147=32'b10111101011001111110001100101001;
	parameter [31:0] W148=32'b10111100010010000001111001110000;
	parameter [31:0] W149=32'b00111010110101000000000101001000;
	parameter [31:0] W150=32'b00111101000111011010111101101100;
	parameter [31:0] W151=32'b00111110011000000111001000110101;
	parameter [31:0] W152=32'b00111101010110110010100111010111;
	parameter [31:0] W153=32'b00111100111001000010010100100011;
	parameter [31:0] W154=32'b00111101101011100110011000100100;
	parameter [31:0] W155=32'b00111101010111100100101011011100;
	parameter [31:0] W156=32'b00111110001000011010100111010000;
	parameter [31:0] W157=32'b00111101110110111010111000001010;
	parameter [31:0] W158=32'b00111101100011100110101001111010;
	parameter [31:0] W159=32'b00111110010001101110111011001001;
	parameter [31:0] W160=32'b00111101100001111011100000010001;
	parameter [31:0] W161=32'b10111100010001010001010101100011;
	parameter [31:0] W162=32'b10111101111110101000110011111100;
	parameter [31:0] W163=32'b10111101101001111101110010000011;
	parameter [31:0] W164=32'b10111110000101011110101000001001;
	parameter [31:0] W165=32'b10111101010101111010000010100111;
	parameter [31:0] W166=32'b10111101011001010101001010100110;
	parameter [31:0] W167=32'b10111101011100110111100111101110;
	parameter [31:0] W168=32'b10111110001000001110011111000010;
	parameter [31:0] W169=32'b00111101001011111111011111001010;
	parameter [31:0] W170=32'b00111101000011011011001110001001;
	parameter [31:0] W171=32'b10111101011101100001001100011011;
	parameter [31:0] W172=32'b10111110100001001010100110110010;
	parameter [31:0] W173=32'b00111100111100011001101110101010;
	parameter [31:0] W174=32'b10111101011111001100111101101000;
	parameter [31:0] W175=32'b10111101110000011001000101000011;
	parameter [31:0] W176=32'b00111100000101101000011000011011;
	parameter [31:0] W177=32'b00111101111001101001101011100011;
	parameter [31:0] W178=32'b00111110100010100000100011011110;
	parameter [31:0] W179=32'b10111011111001110100000011010010;
	parameter [31:0] W180=32'b00111100010101100000111000010101;
	parameter [31:0] W181=32'b00111110010110100010100010010010;
	parameter [31:0] W182=32'b00111111000010111110101010110110;
	parameter [31:0] W183=32'b10111110010011101001100001110000;
	parameter [31:0] W184=32'b10111111001101110000011001011111;
	parameter [31:0] W185=32'b10111111000101001110101100010001;
	parameter [31:0] W186=32'b00111110001000011000000101110101;
	wire [31:0] in0;
	wire [31:0] in1;
	wire [31:0] in2;
	wire [31:0] in3;
	wire [31:0] in4;
	wire [31:0] in5;
	wire [31:0] in6;
	wire [31:0] in7;
	wire [31:0] in8;
	wire [31:0] in9;
	wire [31:0] in10;
	wire [31:0] in11;
	wire [31:0] in12;
	wire [31:0] in13;
	wire [31:0] in14;
	wire [31:0] in15;
	wire [31:0] in16;
	wire [31:0] in17;
	wire [31:0] in18;
	wire [31:0] in19;
	wire [31:0] in20;
	wire [31:0] in21;
	wire [31:0] in22;
	wire [31:0] in23;
	wire [31:0] in24;
	wire [31:0] in25;
	wire [31:0] in26;
	wire [31:0] in27;
	wire [31:0] in28;
	wire [31:0] in29;
	wire [31:0] in30;
	wire [31:0] in31;
	wire [31:0] in32;
	wire [31:0] in33;
	wire [31:0] in34;
	wire [31:0] in35;
	wire [31:0] in36;
	wire [31:0] in37;
	wire [31:0] in38;
	wire [31:0] in39;
	wire [31:0] in40;
	wire [31:0] in41;
	wire [31:0] in42;
	wire [31:0] in43;
	wire [31:0] in44;
	wire [31:0] in45;
	wire [31:0] in46;
	wire [31:0] in47;
	wire [31:0] in48;
	wire [31:0] in49;
	wire [31:0] in50;
	wire [31:0] in51;
	wire [31:0] in52;
	wire [31:0] in53;
	wire [31:0] in54;
	wire [31:0] in55;
	wire [31:0] in56;
	wire [31:0] in57;
	wire [31:0] in58;
	wire [31:0] in59;
	wire [31:0] in60;
	wire [31:0] in61;
	wire [31:0] in62;
	wire [31:0] in63;
	wire [31:0] in64;
	wire [31:0] in65;
	wire [31:0] in66;
	wire [31:0] in67;
	wire [31:0] in68;
	wire [31:0] in69;
	wire [31:0] in70;
	wire [31:0] in71;
	wire [31:0] in72;
	wire [31:0] in73;
	wire [31:0] in74;
	wire [31:0] in75;
	wire [31:0] in76;
	wire [31:0] in77;
	wire [31:0] in78;
	wire [31:0] in79;
	wire [31:0] in80;
	wire [31:0] in81;
	wire [31:0] in82;
	wire [31:0] in83;
	wire [31:0] in84;
	wire [31:0] in85;
	wire [31:0] in86;
	wire [31:0] in87;
	wire [31:0] in88;
	wire [31:0] in89;
	wire [31:0] in90;
	wire [31:0] in91;
	wire [31:0] in92;
	wire [31:0] in93;
	wire [31:0] in94;
	wire [31:0] in95;
	wire [31:0] in96;
	wire [31:0] in97;
	wire [31:0] in98;
	wire [31:0] in99;
	wire [31:0] in100;
	wire [31:0] in101;
	wire [31:0] in102;
	wire [31:0] in103;
	wire [31:0] in104;
	wire [31:0] in105;
	wire [31:0] in106;
	wire [31:0] in107;
	wire [31:0] in108;
	wire [31:0] in109;
	wire [31:0] in110;
	wire [31:0] in111;
	wire [31:0] in112;
	wire [31:0] in113;
	wire [31:0] in114;
	wire [31:0] in115;
	wire [31:0] in116;
	wire [31:0] in117;
	wire [31:0] in118;
	wire [31:0] in119;
	wire [31:0] in120;
	wire [31:0] in121;
	wire [31:0] in122;
	wire [31:0] in123;
	wire [31:0] in124;
	wire [31:0] in125;
	wire [31:0] in126;
	wire [31:0] in127;
	wire [31:0] in128;
	wire [31:0] in129;
	wire [31:0] in130;
	wire [31:0] in131;
	wire [31:0] in132;
	wire [31:0] in133;
	wire [31:0] in134;
	wire [31:0] in135;
	wire [31:0] in136;
	wire [31:0] in137;
	wire [31:0] in138;
	wire [31:0] in139;
	wire [31:0] in140;
	wire [31:0] in141;
	wire [31:0] in142;
	wire [31:0] in143;
	wire [31:0] in144;
	wire [31:0] in145;
	wire [31:0] in146;
	wire [31:0] in147;
	wire [31:0] in148;
	wire [31:0] in149;
	wire [31:0] in150;
	wire [31:0] in151;
	wire [31:0] in152;
	wire [31:0] in153;
	wire [31:0] in154;
	wire [31:0] in155;
	wire [31:0] in156;
	wire [31:0] in157;
	wire [31:0] in158;
	wire [31:0] in159;
	wire [31:0] in160;
	wire [31:0] in161;
	wire [31:0] in162;
	wire [31:0] in163;
	wire [31:0] in164;
	wire [31:0] in165;
	wire [31:0] in166;
	wire [31:0] in167;
	wire [31:0] in168;
	wire [31:0] in169;
	wire [31:0] in170;
	wire [31:0] in171;
	wire [31:0] in172;
	wire [31:0] in173;
	wire [31:0] in174;
	wire [31:0] in175;
	wire [31:0] in176;
	wire [31:0] in177;
	wire [31:0] in178;
	wire [31:0] in179;
	wire [31:0] in180;
	wire [31:0] in181;
	wire [31:0] in182;
	wire [31:0] in183;
	wire [31:0] in184;
	wire [31:0] in185;
	wire [31:0] in186;
	wire [31:0] sum0;
	wire [31:0] sum1;
	wire [31:0] sum2;
	wire [31:0] sum3;
	wire [31:0] sum4;
	wire [31:0] sum5;
	wire [31:0] sum6;
	wire [31:0] sum7;
	wire [31:0] sum8;
	wire [31:0] sum9;
	wire [31:0] sum10;
	wire [31:0] sum11;
	wire [31:0] sum12;
	wire [31:0] sum13;
	wire [31:0] sum14;
	wire [31:0] sum15;
	wire [31:0] sum16;
	wire [31:0] sum17;
	wire [31:0] sum18;
	wire [31:0] sum19;
	wire [31:0] sum20;
	wire [31:0] sum21;
	wire [31:0] sum22;
	wire [31:0] sum23;
	wire [31:0] sum24;
	wire [31:0] sum25;
	wire [31:0] sum26;
	wire [31:0] sum27;
	wire [31:0] sum28;
	wire [31:0] sum29;
	wire [31:0] sum30;
	wire [31:0] sum31;
	wire [31:0] sum32;
	wire [31:0] sum33;
	wire [31:0] sum34;
	wire [31:0] sum35;
	wire [31:0] sum36;
	wire [31:0] sum37;
	wire [31:0] sum38;
	wire [31:0] sum39;
	wire [31:0] sum40;
	wire [31:0] sum41;
	wire [31:0] sum42;
	wire [31:0] sum43;
	wire [31:0] sum44;
	wire [31:0] sum45;
	wire [31:0] sum46;
	wire [31:0] sum47;
	wire [31:0] sum48;
	wire [31:0] sum49;
	wire [31:0] sum50;
	wire [31:0] sum51;
	wire [31:0] sum52;
	wire [31:0] sum53;
	wire [31:0] sum54;
	wire [31:0] sum55;
	wire [31:0] sum56;
	wire [31:0] sum57;
	wire [31:0] sum58;
	wire [31:0] sum59;
	wire [31:0] sum60;
	wire [31:0] sum61;
	wire [31:0] sum62;
	wire [31:0] sum63;
	wire [31:0] sum64;
	wire [31:0] sum65;
	wire [31:0] sum66;
	wire [31:0] sum67;
	wire [31:0] sum68;
	wire [31:0] sum69;
	wire [31:0] sum70;
	wire [31:0] sum71;
	wire [31:0] sum72;
	wire [31:0] sum73;
	wire [31:0] sum74;
	wire [31:0] sum75;
	wire [31:0] sum76;
	wire [31:0] sum77;
	wire [31:0] sum78;
	wire [31:0] sum79;
	wire [31:0] sum80;
	wire [31:0] sum81;
	wire [31:0] sum82;
	wire [31:0] sum83;
	wire [31:0] sum84;
	wire [31:0] sum85;
	wire [31:0] sum86;
	wire [31:0] sum87;
	wire [31:0] sum88;
	wire [31:0] sum89;
	wire [31:0] sum90;
	wire [31:0] sum91;
	wire [31:0] sum92;
	wire [31:0] sum93;
	wire [31:0] sum94;
	wire [31:0] sum95;
	wire [31:0] sum96;
	wire [31:0] sum97;
	wire [31:0] sum98;
	wire [31:0] sum99;
	wire [31:0] sum100;
	wire [31:0] sum101;
	wire [31:0] sum102;
	wire [31:0] sum103;
	wire [31:0] sum104;
	wire [31:0] sum105;
	wire [31:0] sum106;
	wire [31:0] sum107;
	wire [31:0] sum108;
	wire [31:0] sum109;
	wire [31:0] sum110;
	wire [31:0] sum111;
	wire [31:0] sum112;
	wire [31:0] sum113;
	wire [31:0] sum114;
	wire [31:0] sum115;
	wire [31:0] sum116;
	wire [31:0] sum117;
	wire [31:0] sum118;
	wire [31:0] sum119;
	wire [31:0] sum120;
	wire [31:0] sum121;
	wire [31:0] sum122;
	wire [31:0] sum123;
	wire [31:0] sum124;
	wire [31:0] sum125;
	wire [31:0] sum126;
	wire [31:0] sum127;
	wire [31:0] sum128;
	wire [31:0] sum129;
	wire [31:0] sum130;
	wire [31:0] sum131;
	wire [31:0] sum132;
	wire [31:0] sum133;
	wire [31:0] sum134;
	wire [31:0] sum135;
	wire [31:0] sum136;
	wire [31:0] sum137;
	wire [31:0] sum138;
	wire [31:0] sum139;
	wire [31:0] sum140;
	wire [31:0] sum141;
	wire [31:0] sum142;
	wire [31:0] sum143;
	wire [31:0] sum144;
	wire [31:0] sum145;
	wire [31:0] sum146;
	wire [31:0] sum147;
	wire [31:0] sum148;
	wire [31:0] sum149;
	wire [31:0] sum150;
	wire [31:0] sum151;
	wire [31:0] sum152;
	wire [31:0] sum153;
	wire [31:0] sum154;
	wire [31:0] sum155;
	wire [31:0] sum156;
	wire [31:0] sum157;
	wire [31:0] sum158;
	wire [31:0] sum159;
	wire [31:0] sum160;
	wire [31:0] sum161;
	wire [31:0] sum162;
	wire [31:0] sum163;
	wire [31:0] sum164;
	wire [31:0] sum165;
	wire [31:0] sum166;
	wire [31:0] sum167;
	wire [31:0] sum168;
	wire [31:0] sum169;
	wire [31:0] sum170;
	wire [31:0] sum171;
	wire [31:0] sum172;
	wire [31:0] sum173;
	wire [31:0] sum174;
	wire [31:0] sum175;
	wire [31:0] sum176;
	wire [31:0] sum177;
	wire [31:0] sum178;
	wire [31:0] sum179;
	wire [31:0] sum180;
	wire [31:0] sum181;
	wire [31:0] sum182;
	wire [31:0] sum183;
	wire [31:0] sum184;
	wire [31:0] sum185;

	float_mult mult0(
		.x(A0),
		.y(W0),
		.z(in0));
	float_mult mult1(
		.x(A1),
		.y(W1),
		.z(in1));
	float_mult mult2(
		.x(A2),
		.y(W2),
		.z(in2));
	float_mult mult3(
		.x(A3),
		.y(W3),
		.z(in3));
	float_mult mult4(
		.x(A4),
		.y(W4),
		.z(in4));
	float_mult mult5(
		.x(A5),
		.y(W5),
		.z(in5));
	float_mult mult6(
		.x(A6),
		.y(W6),
		.z(in6));
	float_mult mult7(
		.x(A7),
		.y(W7),
		.z(in7));
	float_mult mult8(
		.x(A8),
		.y(W8),
		.z(in8));
	float_mult mult9(
		.x(A9),
		.y(W9),
		.z(in9));
	float_mult mult10(
		.x(A10),
		.y(W10),
		.z(in10));
	float_mult mult11(
		.x(A11),
		.y(W11),
		.z(in11));
	float_mult mult12(
		.x(A12),
		.y(W12),
		.z(in12));
	float_mult mult13(
		.x(A13),
		.y(W13),
		.z(in13));
	float_mult mult14(
		.x(A14),
		.y(W14),
		.z(in14));
	float_mult mult15(
		.x(A15),
		.y(W15),
		.z(in15));
	float_mult mult16(
		.x(A16),
		.y(W16),
		.z(in16));
	float_mult mult17(
		.x(A17),
		.y(W17),
		.z(in17));
	float_mult mult18(
		.x(A18),
		.y(W18),
		.z(in18));
	float_mult mult19(
		.x(A19),
		.y(W19),
		.z(in19));
	float_mult mult20(
		.x(A20),
		.y(W20),
		.z(in20));
	float_mult mult21(
		.x(A21),
		.y(W21),
		.z(in21));
	float_mult mult22(
		.x(A22),
		.y(W22),
		.z(in22));
	float_mult mult23(
		.x(A23),
		.y(W23),
		.z(in23));
	float_mult mult24(
		.x(A24),
		.y(W24),
		.z(in24));
	float_mult mult25(
		.x(A25),
		.y(W25),
		.z(in25));
	float_mult mult26(
		.x(A26),
		.y(W26),
		.z(in26));
	float_mult mult27(
		.x(A27),
		.y(W27),
		.z(in27));
	float_mult mult28(
		.x(A28),
		.y(W28),
		.z(in28));
	float_mult mult29(
		.x(A29),
		.y(W29),
		.z(in29));
	float_mult mult30(
		.x(A30),
		.y(W30),
		.z(in30));
	float_mult mult31(
		.x(A31),
		.y(W31),
		.z(in31));
	float_mult mult32(
		.x(A32),
		.y(W32),
		.z(in32));
	float_mult mult33(
		.x(A33),
		.y(W33),
		.z(in33));
	float_mult mult34(
		.x(A34),
		.y(W34),
		.z(in34));
	float_mult mult35(
		.x(A35),
		.y(W35),
		.z(in35));
	float_mult mult36(
		.x(A36),
		.y(W36),
		.z(in36));
	float_mult mult37(
		.x(A37),
		.y(W37),
		.z(in37));
	float_mult mult38(
		.x(A38),
		.y(W38),
		.z(in38));
	float_mult mult39(
		.x(A39),
		.y(W39),
		.z(in39));
	float_mult mult40(
		.x(A40),
		.y(W40),
		.z(in40));
	float_mult mult41(
		.x(A41),
		.y(W41),
		.z(in41));
	float_mult mult42(
		.x(A42),
		.y(W42),
		.z(in42));
	float_mult mult43(
		.x(A43),
		.y(W43),
		.z(in43));
	float_mult mult44(
		.x(A44),
		.y(W44),
		.z(in44));
	float_mult mult45(
		.x(A45),
		.y(W45),
		.z(in45));
	float_mult mult46(
		.x(A46),
		.y(W46),
		.z(in46));
	float_mult mult47(
		.x(A47),
		.y(W47),
		.z(in47));
	float_mult mult48(
		.x(A48),
		.y(W48),
		.z(in48));
	float_mult mult49(
		.x(A49),
		.y(W49),
		.z(in49));
	float_mult mult50(
		.x(A50),
		.y(W50),
		.z(in50));
	float_mult mult51(
		.x(A51),
		.y(W51),
		.z(in51));
	float_mult mult52(
		.x(A52),
		.y(W52),
		.z(in52));
	float_mult mult53(
		.x(A53),
		.y(W53),
		.z(in53));
	float_mult mult54(
		.x(A54),
		.y(W54),
		.z(in54));
	float_mult mult55(
		.x(A55),
		.y(W55),
		.z(in55));
	float_mult mult56(
		.x(A56),
		.y(W56),
		.z(in56));
	float_mult mult57(
		.x(A57),
		.y(W57),
		.z(in57));
	float_mult mult58(
		.x(A58),
		.y(W58),
		.z(in58));
	float_mult mult59(
		.x(A59),
		.y(W59),
		.z(in59));
	float_mult mult60(
		.x(A60),
		.y(W60),
		.z(in60));
	float_mult mult61(
		.x(A61),
		.y(W61),
		.z(in61));
	float_mult mult62(
		.x(A62),
		.y(W62),
		.z(in62));
	float_mult mult63(
		.x(A63),
		.y(W63),
		.z(in63));
	float_mult mult64(
		.x(A64),
		.y(W64),
		.z(in64));
	float_mult mult65(
		.x(A65),
		.y(W65),
		.z(in65));
	float_mult mult66(
		.x(A66),
		.y(W66),
		.z(in66));
	float_mult mult67(
		.x(A67),
		.y(W67),
		.z(in67));
	float_mult mult68(
		.x(A68),
		.y(W68),
		.z(in68));
	float_mult mult69(
		.x(A69),
		.y(W69),
		.z(in69));
	float_mult mult70(
		.x(A70),
		.y(W70),
		.z(in70));
	float_mult mult71(
		.x(A71),
		.y(W71),
		.z(in71));
	float_mult mult72(
		.x(A72),
		.y(W72),
		.z(in72));
	float_mult mult73(
		.x(A73),
		.y(W73),
		.z(in73));
	float_mult mult74(
		.x(A74),
		.y(W74),
		.z(in74));
	float_mult mult75(
		.x(A75),
		.y(W75),
		.z(in75));
	float_mult mult76(
		.x(A76),
		.y(W76),
		.z(in76));
	float_mult mult77(
		.x(A77),
		.y(W77),
		.z(in77));
	float_mult mult78(
		.x(A78),
		.y(W78),
		.z(in78));
	float_mult mult79(
		.x(A79),
		.y(W79),
		.z(in79));
	float_mult mult80(
		.x(A80),
		.y(W80),
		.z(in80));
	float_mult mult81(
		.x(A81),
		.y(W81),
		.z(in81));
	float_mult mult82(
		.x(A82),
		.y(W82),
		.z(in82));
	float_mult mult83(
		.x(A83),
		.y(W83),
		.z(in83));
	float_mult mult84(
		.x(A84),
		.y(W84),
		.z(in84));
	float_mult mult85(
		.x(A85),
		.y(W85),
		.z(in85));
	float_mult mult86(
		.x(A86),
		.y(W86),
		.z(in86));
	float_mult mult87(
		.x(A87),
		.y(W87),
		.z(in87));
	float_mult mult88(
		.x(A88),
		.y(W88),
		.z(in88));
	float_mult mult89(
		.x(A89),
		.y(W89),
		.z(in89));
	float_mult mult90(
		.x(A90),
		.y(W90),
		.z(in90));
	float_mult mult91(
		.x(A91),
		.y(W91),
		.z(in91));
	float_mult mult92(
		.x(A92),
		.y(W92),
		.z(in92));
	float_mult mult93(
		.x(A93),
		.y(W93),
		.z(in93));
	float_mult mult94(
		.x(A94),
		.y(W94),
		.z(in94));
	float_mult mult95(
		.x(A95),
		.y(W95),
		.z(in95));
	float_mult mult96(
		.x(A96),
		.y(W96),
		.z(in96));
	float_mult mult97(
		.x(A97),
		.y(W97),
		.z(in97));
	float_mult mult98(
		.x(A98),
		.y(W98),
		.z(in98));
	float_mult mult99(
		.x(A99),
		.y(W99),
		.z(in99));
	float_mult mult100(
		.x(A100),
		.y(W100),
		.z(in100));
	float_mult mult101(
		.x(A101),
		.y(W101),
		.z(in101));
	float_mult mult102(
		.x(A102),
		.y(W102),
		.z(in102));
	float_mult mult103(
		.x(A103),
		.y(W103),
		.z(in103));
	float_mult mult104(
		.x(A104),
		.y(W104),
		.z(in104));
	float_mult mult105(
		.x(A105),
		.y(W105),
		.z(in105));
	float_mult mult106(
		.x(A106),
		.y(W106),
		.z(in106));
	float_mult mult107(
		.x(A107),
		.y(W107),
		.z(in107));
	float_mult mult108(
		.x(A108),
		.y(W108),
		.z(in108));
	float_mult mult109(
		.x(A109),
		.y(W109),
		.z(in109));
	float_mult mult110(
		.x(A110),
		.y(W110),
		.z(in110));
	float_mult mult111(
		.x(A111),
		.y(W111),
		.z(in111));
	float_mult mult112(
		.x(A112),
		.y(W112),
		.z(in112));
	float_mult mult113(
		.x(A113),
		.y(W113),
		.z(in113));
	float_mult mult114(
		.x(A114),
		.y(W114),
		.z(in114));
	float_mult mult115(
		.x(A115),
		.y(W115),
		.z(in115));
	float_mult mult116(
		.x(A116),
		.y(W116),
		.z(in116));
	float_mult mult117(
		.x(A117),
		.y(W117),
		.z(in117));
	float_mult mult118(
		.x(A118),
		.y(W118),
		.z(in118));
	float_mult mult119(
		.x(A119),
		.y(W119),
		.z(in119));
	float_mult mult120(
		.x(A120),
		.y(W120),
		.z(in120));
	float_mult mult121(
		.x(A121),
		.y(W121),
		.z(in121));
	float_mult mult122(
		.x(A122),
		.y(W122),
		.z(in122));
	float_mult mult123(
		.x(A123),
		.y(W123),
		.z(in123));
	float_mult mult124(
		.x(A124),
		.y(W124),
		.z(in124));
	float_mult mult125(
		.x(A125),
		.y(W125),
		.z(in125));
	float_mult mult126(
		.x(A126),
		.y(W126),
		.z(in126));
	float_mult mult127(
		.x(A127),
		.y(W127),
		.z(in127));
	float_mult mult128(
		.x(A128),
		.y(W128),
		.z(in128));
	float_mult mult129(
		.x(A129),
		.y(W129),
		.z(in129));
	float_mult mult130(
		.x(A130),
		.y(W130),
		.z(in130));
	float_mult mult131(
		.x(A131),
		.y(W131),
		.z(in131));
	float_mult mult132(
		.x(A132),
		.y(W132),
		.z(in132));
	float_mult mult133(
		.x(A133),
		.y(W133),
		.z(in133));
	float_mult mult134(
		.x(A134),
		.y(W134),
		.z(in134));
	float_mult mult135(
		.x(A135),
		.y(W135),
		.z(in135));
	float_mult mult136(
		.x(A136),
		.y(W136),
		.z(in136));
	float_mult mult137(
		.x(A137),
		.y(W137),
		.z(in137));
	float_mult mult138(
		.x(A138),
		.y(W138),
		.z(in138));
	float_mult mult139(
		.x(A139),
		.y(W139),
		.z(in139));
	float_mult mult140(
		.x(A140),
		.y(W140),
		.z(in140));
	float_mult mult141(
		.x(A141),
		.y(W141),
		.z(in141));
	float_mult mult142(
		.x(A142),
		.y(W142),
		.z(in142));
	float_mult mult143(
		.x(A143),
		.y(W143),
		.z(in143));
	float_mult mult144(
		.x(A144),
		.y(W144),
		.z(in144));
	float_mult mult145(
		.x(A145),
		.y(W145),
		.z(in145));
	float_mult mult146(
		.x(A146),
		.y(W146),
		.z(in146));
	float_mult mult147(
		.x(A147),
		.y(W147),
		.z(in147));
	float_mult mult148(
		.x(A148),
		.y(W148),
		.z(in148));
	float_mult mult149(
		.x(A149),
		.y(W149),
		.z(in149));
	float_mult mult150(
		.x(A150),
		.y(W150),
		.z(in150));
	float_mult mult151(
		.x(A151),
		.y(W151),
		.z(in151));
	float_mult mult152(
		.x(A152),
		.y(W152),
		.z(in152));
	float_mult mult153(
		.x(A153),
		.y(W153),
		.z(in153));
	float_mult mult154(
		.x(A154),
		.y(W154),
		.z(in154));
	float_mult mult155(
		.x(A155),
		.y(W155),
		.z(in155));
	float_mult mult156(
		.x(A156),
		.y(W156),
		.z(in156));
	float_mult mult157(
		.x(A157),
		.y(W157),
		.z(in157));
	float_mult mult158(
		.x(A158),
		.y(W158),
		.z(in158));
	float_mult mult159(
		.x(A159),
		.y(W159),
		.z(in159));
	float_mult mult160(
		.x(A160),
		.y(W160),
		.z(in160));
	float_mult mult161(
		.x(A161),
		.y(W161),
		.z(in161));
	float_mult mult162(
		.x(A162),
		.y(W162),
		.z(in162));
	float_mult mult163(
		.x(A163),
		.y(W163),
		.z(in163));
	float_mult mult164(
		.x(A164),
		.y(W164),
		.z(in164));
	float_mult mult165(
		.x(A165),
		.y(W165),
		.z(in165));
	float_mult mult166(
		.x(A166),
		.y(W166),
		.z(in166));
	float_mult mult167(
		.x(A167),
		.y(W167),
		.z(in167));
	float_mult mult168(
		.x(A168),
		.y(W168),
		.z(in168));
	float_mult mult169(
		.x(A169),
		.y(W169),
		.z(in169));
	float_mult mult170(
		.x(A170),
		.y(W170),
		.z(in170));
	float_mult mult171(
		.x(A171),
		.y(W171),
		.z(in171));
	float_mult mult172(
		.x(A172),
		.y(W172),
		.z(in172));
	float_mult mult173(
		.x(A173),
		.y(W173),
		.z(in173));
	float_mult mult174(
		.x(A174),
		.y(W174),
		.z(in174));
	float_mult mult175(
		.x(A175),
		.y(W175),
		.z(in175));
	float_mult mult176(
		.x(A176),
		.y(W176),
		.z(in176));
	float_mult mult177(
		.x(A177),
		.y(W177),
		.z(in177));
	float_mult mult178(
		.x(A178),
		.y(W178),
		.z(in178));
	float_mult mult179(
		.x(A179),
		.y(W179),
		.z(in179));
	float_mult mult180(
		.x(A180),
		.y(W180),
		.z(in180));
	float_mult mult181(
		.x(A181),
		.y(W181),
		.z(in181));
	float_mult mult182(
		.x(A182),
		.y(W182),
		.z(in182));
	float_mult mult183(
		.x(A183),
		.y(W183),
		.z(in183));
	float_mult mult184(
		.x(A184),
		.y(W184),
		.z(in184));
	float_mult mult185(
		.x(A185),
		.y(W185),
		.z(in185));
	float_mult mult186(
		.x(A186),
		.y(W186),
		.z(in186));

	float_adder add0(
		.a(in0),
		.b(in1),
		.Out(sum0),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add1(
		.a(in2),
		.b(in3),
		.Out(sum1),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add2(
		.a(in4),
		.b(in5),
		.Out(sum2),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add3(
		.a(in6),
		.b(in7),
		.Out(sum3),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add4(
		.a(in8),
		.b(in9),
		.Out(sum4),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add5(
		.a(in10),
		.b(in11),
		.Out(sum5),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add6(
		.a(in12),
		.b(in13),
		.Out(sum6),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add7(
		.a(in14),
		.b(in15),
		.Out(sum7),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add8(
		.a(in16),
		.b(in17),
		.Out(sum8),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add9(
		.a(in18),
		.b(in19),
		.Out(sum9),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add10(
		.a(in20),
		.b(in21),
		.Out(sum10),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add11(
		.a(in22),
		.b(in23),
		.Out(sum11),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add12(
		.a(in24),
		.b(in25),
		.Out(sum12),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add13(
		.a(in26),
		.b(in27),
		.Out(sum13),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add14(
		.a(in28),
		.b(in29),
		.Out(sum14),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add15(
		.a(in30),
		.b(in31),
		.Out(sum15),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add16(
		.a(in32),
		.b(in33),
		.Out(sum16),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add17(
		.a(in34),
		.b(in35),
		.Out(sum17),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add18(
		.a(in36),
		.b(in37),
		.Out(sum18),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add19(
		.a(in38),
		.b(in39),
		.Out(sum19),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add20(
		.a(in40),
		.b(in41),
		.Out(sum20),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add21(
		.a(in42),
		.b(in43),
		.Out(sum21),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add22(
		.a(in44),
		.b(in45),
		.Out(sum22),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add23(
		.a(in46),
		.b(in47),
		.Out(sum23),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add24(
		.a(in48),
		.b(in49),
		.Out(sum24),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add25(
		.a(in50),
		.b(in51),
		.Out(sum25),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add26(
		.a(in52),
		.b(in53),
		.Out(sum26),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add27(
		.a(in54),
		.b(in55),
		.Out(sum27),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add28(
		.a(in56),
		.b(in57),
		.Out(sum28),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add29(
		.a(in58),
		.b(in59),
		.Out(sum29),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add30(
		.a(in60),
		.b(in61),
		.Out(sum30),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add31(
		.a(in62),
		.b(in63),
		.Out(sum31),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add32(
		.a(in64),
		.b(in65),
		.Out(sum32),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add33(
		.a(in66),
		.b(in67),
		.Out(sum33),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add34(
		.a(in68),
		.b(in69),
		.Out(sum34),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add35(
		.a(in70),
		.b(in71),
		.Out(sum35),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add36(
		.a(in72),
		.b(in73),
		.Out(sum36),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add37(
		.a(in74),
		.b(in75),
		.Out(sum37),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add38(
		.a(in76),
		.b(in77),
		.Out(sum38),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add39(
		.a(in78),
		.b(in79),
		.Out(sum39),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add40(
		.a(in80),
		.b(in81),
		.Out(sum40),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add41(
		.a(in82),
		.b(in83),
		.Out(sum41),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add42(
		.a(in84),
		.b(in85),
		.Out(sum42),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add43(
		.a(in86),
		.b(in87),
		.Out(sum43),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add44(
		.a(in88),
		.b(in89),
		.Out(sum44),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add45(
		.a(in90),
		.b(in91),
		.Out(sum45),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add46(
		.a(in92),
		.b(in93),
		.Out(sum46),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add47(
		.a(in94),
		.b(in95),
		.Out(sum47),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add48(
		.a(in96),
		.b(in97),
		.Out(sum48),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add49(
		.a(in98),
		.b(in99),
		.Out(sum49),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add50(
		.a(in100),
		.b(in101),
		.Out(sum50),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add51(
		.a(in102),
		.b(in103),
		.Out(sum51),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add52(
		.a(in104),
		.b(in105),
		.Out(sum52),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add53(
		.a(in106),
		.b(in107),
		.Out(sum53),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add54(
		.a(in108),
		.b(in109),
		.Out(sum54),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add55(
		.a(in110),
		.b(in111),
		.Out(sum55),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add56(
		.a(in112),
		.b(in113),
		.Out(sum56),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add57(
		.a(in114),
		.b(in115),
		.Out(sum57),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add58(
		.a(in116),
		.b(in117),
		.Out(sum58),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add59(
		.a(in118),
		.b(in119),
		.Out(sum59),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add60(
		.a(in120),
		.b(in121),
		.Out(sum60),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add61(
		.a(in122),
		.b(in123),
		.Out(sum61),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add62(
		.a(in124),
		.b(in125),
		.Out(sum62),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add63(
		.a(in126),
		.b(in127),
		.Out(sum63),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add64(
		.a(in128),
		.b(in129),
		.Out(sum64),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add65(
		.a(in130),
		.b(in131),
		.Out(sum65),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add66(
		.a(in132),
		.b(in133),
		.Out(sum66),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add67(
		.a(in134),
		.b(in135),
		.Out(sum67),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add68(
		.a(in136),
		.b(in137),
		.Out(sum68),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add69(
		.a(in138),
		.b(in139),
		.Out(sum69),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add70(
		.a(in140),
		.b(in141),
		.Out(sum70),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add71(
		.a(in142),
		.b(in143),
		.Out(sum71),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add72(
		.a(in144),
		.b(in145),
		.Out(sum72),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add73(
		.a(in146),
		.b(in147),
		.Out(sum73),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add74(
		.a(in148),
		.b(in149),
		.Out(sum74),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add75(
		.a(in150),
		.b(in151),
		.Out(sum75),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add76(
		.a(in152),
		.b(in153),
		.Out(sum76),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add77(
		.a(in154),
		.b(in155),
		.Out(sum77),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add78(
		.a(in156),
		.b(in157),
		.Out(sum78),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add79(
		.a(in158),
		.b(in159),
		.Out(sum79),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add80(
		.a(in160),
		.b(in161),
		.Out(sum80),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add81(
		.a(in162),
		.b(in163),
		.Out(sum81),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add82(
		.a(in164),
		.b(in165),
		.Out(sum82),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add83(
		.a(in166),
		.b(in167),
		.Out(sum83),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add84(
		.a(in168),
		.b(in169),
		.Out(sum84),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add85(
		.a(in170),
		.b(in171),
		.Out(sum85),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add86(
		.a(in172),
		.b(in173),
		.Out(sum86),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add87(
		.a(in174),
		.b(in175),
		.Out(sum87),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add88(
		.a(in176),
		.b(in177),
		.Out(sum88),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add89(
		.a(in178),
		.b(in179),
		.Out(sum89),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add90(
		.a(in180),
		.b(in181),
		.Out(sum90),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add91(
		.a(in182),
		.b(in183),
		.Out(sum91),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add92(
		.a(in184),
		.b(in185),
		.Out(sum92),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add93(
		.a(sum0),
		.b(sum1),
		.Out(sum93),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add94(
		.a(sum2),
		.b(sum3),
		.Out(sum94),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add95(
		.a(sum4),
		.b(sum5),
		.Out(sum95),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add96(
		.a(sum6),
		.b(sum7),
		.Out(sum96),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add97(
		.a(sum8),
		.b(sum9),
		.Out(sum97),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add98(
		.a(sum10),
		.b(sum11),
		.Out(sum98),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add99(
		.a(sum12),
		.b(sum13),
		.Out(sum99),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add100(
		.a(sum14),
		.b(sum15),
		.Out(sum100),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add101(
		.a(sum16),
		.b(sum17),
		.Out(sum101),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add102(
		.a(sum18),
		.b(sum19),
		.Out(sum102),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add103(
		.a(sum20),
		.b(sum21),
		.Out(sum103),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add104(
		.a(sum22),
		.b(sum23),
		.Out(sum104),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add105(
		.a(sum24),
		.b(sum25),
		.Out(sum105),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add106(
		.a(sum26),
		.b(sum27),
		.Out(sum106),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add107(
		.a(sum28),
		.b(sum29),
		.Out(sum107),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add108(
		.a(sum30),
		.b(sum31),
		.Out(sum108),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add109(
		.a(sum32),
		.b(sum33),
		.Out(sum109),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add110(
		.a(sum34),
		.b(sum35),
		.Out(sum110),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add111(
		.a(sum36),
		.b(sum37),
		.Out(sum111),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add112(
		.a(sum38),
		.b(sum39),
		.Out(sum112),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add113(
		.a(sum40),
		.b(sum41),
		.Out(sum113),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add114(
		.a(sum42),
		.b(sum43),
		.Out(sum114),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add115(
		.a(sum44),
		.b(sum45),
		.Out(sum115),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add116(
		.a(sum46),
		.b(sum47),
		.Out(sum116),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add117(
		.a(sum48),
		.b(sum49),
		.Out(sum117),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add118(
		.a(sum50),
		.b(sum51),
		.Out(sum118),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add119(
		.a(sum52),
		.b(sum53),
		.Out(sum119),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add120(
		.a(sum54),
		.b(sum55),
		.Out(sum120),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add121(
		.a(sum56),
		.b(sum57),
		.Out(sum121),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add122(
		.a(sum58),
		.b(sum59),
		.Out(sum122),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add123(
		.a(sum60),
		.b(sum61),
		.Out(sum123),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add124(
		.a(sum62),
		.b(sum63),
		.Out(sum124),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add125(
		.a(sum64),
		.b(sum65),
		.Out(sum125),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add126(
		.a(sum66),
		.b(sum67),
		.Out(sum126),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add127(
		.a(sum68),
		.b(sum69),
		.Out(sum127),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add128(
		.a(sum70),
		.b(sum71),
		.Out(sum128),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add129(
		.a(sum72),
		.b(sum73),
		.Out(sum129),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add130(
		.a(sum74),
		.b(sum75),
		.Out(sum130),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add131(
		.a(sum76),
		.b(sum77),
		.Out(sum131),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add132(
		.a(sum78),
		.b(sum79),
		.Out(sum132),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add133(
		.a(sum80),
		.b(sum81),
		.Out(sum133),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add134(
		.a(sum82),
		.b(sum83),
		.Out(sum134),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add135(
		.a(sum84),
		.b(sum85),
		.Out(sum135),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add136(
		.a(sum86),
		.b(sum87),
		.Out(sum136),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add137(
		.a(sum88),
		.b(sum89),
		.Out(sum137),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add138(
		.a(sum90),
		.b(sum91),
		.Out(sum138),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add139(
		.a(sum92),
		.b(in186),
		.Out(sum139),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add140(
		.a(sum93),
		.b(sum94),
		.Out(sum140),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add141(
		.a(sum95),
		.b(sum96),
		.Out(sum141),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add142(
		.a(sum97),
		.b(sum98),
		.Out(sum142),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add143(
		.a(sum99),
		.b(sum100),
		.Out(sum143),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add144(
		.a(sum101),
		.b(sum102),
		.Out(sum144),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add145(
		.a(sum103),
		.b(sum104),
		.Out(sum145),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add146(
		.a(sum105),
		.b(sum106),
		.Out(sum146),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add147(
		.a(sum107),
		.b(sum108),
		.Out(sum147),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add148(
		.a(sum109),
		.b(sum110),
		.Out(sum148),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add149(
		.a(sum111),
		.b(sum112),
		.Out(sum149),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add150(
		.a(sum113),
		.b(sum114),
		.Out(sum150),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add151(
		.a(sum115),
		.b(sum116),
		.Out(sum151),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add152(
		.a(sum117),
		.b(sum118),
		.Out(sum152),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add153(
		.a(sum119),
		.b(sum120),
		.Out(sum153),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add154(
		.a(sum121),
		.b(sum122),
		.Out(sum154),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add155(
		.a(sum123),
		.b(sum124),
		.Out(sum155),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add156(
		.a(sum125),
		.b(sum126),
		.Out(sum156),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add157(
		.a(sum127),
		.b(sum128),
		.Out(sum157),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add158(
		.a(sum129),
		.b(sum130),
		.Out(sum158),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add159(
		.a(sum131),
		.b(sum132),
		.Out(sum159),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add160(
		.a(sum133),
		.b(sum134),
		.Out(sum160),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add161(
		.a(sum135),
		.b(sum136),
		.Out(sum161),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add162(
		.a(sum137),
		.b(sum138),
		.Out(sum162),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add163(
		.a(sum140),
		.b(sum141),
		.Out(sum163),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add164(
		.a(sum142),
		.b(sum143),
		.Out(sum164),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add165(
		.a(sum144),
		.b(sum145),
		.Out(sum165),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add166(
		.a(sum146),
		.b(sum147),
		.Out(sum166),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add167(
		.a(sum148),
		.b(sum149),
		.Out(sum167),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add168(
		.a(sum150),
		.b(sum151),
		.Out(sum168),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add169(
		.a(sum152),
		.b(sum153),
		.Out(sum169),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add170(
		.a(sum154),
		.b(sum155),
		.Out(sum170),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add171(
		.a(sum156),
		.b(sum157),
		.Out(sum171),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add172(
		.a(sum158),
		.b(sum159),
		.Out(sum172),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add173(
		.a(sum160),
		.b(sum161),
		.Out(sum173),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add174(
		.a(sum162),
		.b(sum139),
		.Out(sum174),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add175(
		.a(sum163),
		.b(sum164),
		.Out(sum175),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add176(
		.a(sum165),
		.b(sum166),
		.Out(sum176),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add177(
		.a(sum167),
		.b(sum168),
		.Out(sum177),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add178(
		.a(sum169),
		.b(sum170),
		.Out(sum178),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add179(
		.a(sum171),
		.b(sum172),
		.Out(sum179),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add180(
		.a(sum173),
		.b(sum174),
		.Out(sum180),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add181(
		.a(sum175),
		.b(sum176),
		.Out(sum181),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add182(
		.a(sum177),
		.b(sum178),
		.Out(sum182),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add183(
		.a(sum179),
		.b(sum180),
		.Out(sum183),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add184(
		.a(sum181),
		.b(sum182),
		.Out(sum184),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add185(
		.a(sum184),
		.b(sum183),
		.Out(N1),
		.Out_test(),
		.shift(),
		.c_out());
always@(*)
	begin 
		if(N1[31]==0)
			N1=N1;
		else
			N1=32'd0;
	end
endmodule
