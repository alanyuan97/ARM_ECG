module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 4097;
	I1x = -7625;
	I2x = 3158;
	I3x = -7382;
	I4x = 4859;
	I5x = -4745;
	I6x = 1257;
	I7x = 6516;
	I8x = -306;
	I9x = -2935;
	I10x = -7870;
	I11x = -2682;
	I12x = -1913;
	I13x = -4451;
	I14x = -2907;
	I15x = -6335;
	I16x = -4923;
	I17x = 4684;
	I18x = -2293;
	I19x = 1603;
	I20x = 7672;
	I21x = 522;
	I22x = -4544;
	I23x = -5713;
	I24x = -911;
	I25x = 6274;
	I26x = 2285;
	I27x = -1714;
	I28x = 3605;
	I29x = 7202;
	I30x = -6591;
	I31x = -5532;
	I32x = -3374;
	I33x = -2596;
	I34x = 4078;
	I35x = 5436;
	I36x = -7492;
	I37x = 2241;
	I38x = 6369;
	I39x = 4653;
	I40x = 5715;
	I41x = -5142;
	I42x = -2939;
	I43x = 3596;
	I44x = 5506;
	I45x = -1224;
	I46x = -7803;
	I47x = 997;
	I48x = -4566;
	I49x = -561;
	I50x = 7895;
	I51x = -1649;
	I52x = -7105;
	I53x = -7523;
	I54x = 5648;
	I55x = 1851;
	I56x = 2937;
	I57x = 4086;
	I58x = -7623;
	I59x = -5570;
	I60x = 2735;
	I61x = 5682;
	I62x = -5085;
	I63x = -4487;
	I64x = -3125;
	I65x = 3109;
	I66x = -5252;
	I67x = -3692;
	I68x = -6364;
	I69x = 4675;
	I70x = -5566;
	I71x = 3783;
	I72x = -3742;
	I73x = -2481;
	I74x = 2545;
	I75x = -6518;
	I76x = -6026;
	I77x = 5782;
	I78x = -1085;
	I79x = 4511;
	I80x = 1739;
	I81x = -6916;
	I82x = -4082;
	I83x = 350;
	I84x = 85;
	I85x = -5322;
	I86x = 7592;
	I87x = -4362;
	I88x = 5517;
	I89x = 3541;
	I90x = -2729;
	I91x = -2834;
	I92x = 7040;
	I93x = -560;
	I94x = 6802;
	I95x = -5741;
	I96x = 169;
	I97x = 5987;
	I98x = -2485;
	I99x = -3931;
	I100x = -3706;
	I101x = 7085;
	I102x = -6085;
	I103x = 7058;
	I104x = 771;
	I105x = -6231;
	I106x = 390;
	I107x = 114;
	I108x = 4018;
	I109x = 6650;
	I110x = 7450;
	I111x = 6049;
	I112x = -2971;
	I113x = 4139;
	I114x = -6664;
	I115x = -1155;
	I116x = -494;
	I117x = -7121;
	I118x = -7464;
	I119x = -2829;
	I120x = -4939;
	I121x = 5547;
	I122x = 3551;
	I123x = 230;
	I124x = -5708;
	I125x = -3046;
	I126x = -3523;
	I127x = -6494;
	I128x = 6154;
	I129x = 7491;
	I130x = -5873;
	I131x = -5120;
	I132x = -6381;
	I133x = -889;
	I134x = 2201;
	I135x = 2794;
	I136x = 4632;
	I137x = -6042;
	I138x = -1372;
	I139x = 3393;
	I140x = -2318;
	I141x = -223;
	I142x = -1900;
	I143x = 6452;
	I144x = 6070;
	I145x = 2471;
	I146x = 2797;
	I147x = -7191;
	I148x = -2129;
	I149x = 6794;
	I150x = -7649;
	I151x = 2879;
	I152x = 2085;
	I153x = -6913;
	I154x = 4665;
	I155x = -4450;
	I156x = 7289;
	I157x = -6375;
	I158x = -2988;
	I159x = 5065;
	I160x = -5044;
	I161x = 2143;
	I162x = -1213;
	I163x = 3940;
	I164x = 6879;
	I165x = -8085;
	I166x = 2039;
	I167x = 2835;
	I168x = -5052;
	I169x = -4640;
	I170x = 6925;
	I171x = 4700;
	I172x = -2320;
	I173x = -5883;
	I174x = -5660;
	I175x = 1619;
	I176x = 7948;
	I177x = 1957;
	I178x = 3563;
	I179x = -6344;
	I180x = -5555;
	I181x = -5967;
	I182x = 6847;
	I183x = -3155;
	I184x = 2313;
	I185x = -2091;
	I186x = -7251;
	end
endmodule
[0.        0.        0.2413817 0.        0.       ] 

 [0, 0, 1977, 0, 0] 

 ['0000000000000000', '0000000000000000', '0000011110111001', '0000000000000000', '0000000000000000']
