module node1_1(clk,N1x,A0x,A1x,A2x,A3x,A4x,A5x,A6x,A7x,A8x,A9x,A10x,A11x,A12x,A13x,A14x,A15x,A16x,A17x,A18x,A19x,A20x,A21x,A22x,A23x,A24x,A25x,A26x,A27x,A28x,A29x,A30x,A31x,A32x,A33x,A34x,A35x,A36x,A37x,A38x,A39x,A40x,A41x,A42x,A43x,A44x,A45x,A46x,A47x,A48x,A49x,A50x,A51x,A52x,A53x,A54x,A55x,A56x,A57x,A58x,A59x,A60x,A61x,A62x,A63x,A64x,A65x,A66x,A67x,A68x,A69x,A70x,A71x,A72x,A73x,A74x,A75x,A76x,A77x,A78x,A79x,A80x,A81x,A82x,A83x,A84x,A85x,A86x,A87x,A88x,A89x,A90x,A91x,A92x,A93x,A94x,A95x,A96x,A97x,A98x,A99x,A100x,A101x,A102x,A103x,A104x,A105x,A106x,A107x,A108x,A109x,A110x,A111x,A112x,A113x,A114x,A115x,A116x,A117x,A118x,A119x,A120x,A121x,A122x,A123x,A124x,A125x,A126x,A127x,A128x,A129x,A130x,A131x,A132x,A133x,A134x,A135x,A136x,A137x,A138x,A139x,A140x,A141x,A142x,A143x,A144x,A145x,A146x,A147x,A148x,A149x,A150x,A151x,A152x,A153x,A154x,A155x,A156x,A157x,A158x,A159x,A160x,A161x,A162x,A163x,A164x,A165x,A166x,A167x,A168x,A169x,A170x,A171x,A172x,A173x,A174x,A175x,A176x,A177x,A178x,A179x,A180x,A181x,A182x,A183x,A184x,A185x,A186x);
	input clk;
	input [31:0] A0x;
	input clk;
	input [31:0] A1x;
	input clk;
	input [31:0] A2x;
	input clk;
	input [31:0] A3x;
	input clk;
	input [31:0] A4x;
	input clk;
	input [31:0] A5x;
	input clk;
	input [31:0] A6x;
	input clk;
	input [31:0] A7x;
	input clk;
	input [31:0] A8x;
	input clk;
	input [31:0] A9x;
	input clk;
	input [31:0] A10x;
	input clk;
	input [31:0] A11x;
	input clk;
	input [31:0] A12x;
	input clk;
	input [31:0] A13x;
	input clk;
	input [31:0] A14x;
	input clk;
	input [31:0] A15x;
	input clk;
	input [31:0] A16x;
	input clk;
	input [31:0] A17x;
	input clk;
	input [31:0] A18x;
	input clk;
	input [31:0] A19x;
	input clk;
	input [31:0] A20x;
	input clk;
	input [31:0] A21x;
	input clk;
	input [31:0] A22x;
	input clk;
	input [31:0] A23x;
	input clk;
	input [31:0] A24x;
	input clk;
	input [31:0] A25x;
	input clk;
	input [31:0] A26x;
	input clk;
	input [31:0] A27x;
	input clk;
	input [31:0] A28x;
	input clk;
	input [31:0] A29x;
	input clk;
	input [31:0] A30x;
	input clk;
	input [31:0] A31x;
	input clk;
	input [31:0] A32x;
	input clk;
	input [31:0] A33x;
	input clk;
	input [31:0] A34x;
	input clk;
	input [31:0] A35x;
	input clk;
	input [31:0] A36x;
	input clk;
	input [31:0] A37x;
	input clk;
	input [31:0] A38x;
	input clk;
	input [31:0] A39x;
	input clk;
	input [31:0] A40x;
	input clk;
	input [31:0] A41x;
	input clk;
	input [31:0] A42x;
	input clk;
	input [31:0] A43x;
	input clk;
	input [31:0] A44x;
	input clk;
	input [31:0] A45x;
	input clk;
	input [31:0] A46x;
	input clk;
	input [31:0] A47x;
	input clk;
	input [31:0] A48x;
	input clk;
	input [31:0] A49x;
	input clk;
	input [31:0] A50x;
	input clk;
	input [31:0] A51x;
	input clk;
	input [31:0] A52x;
	input clk;
	input [31:0] A53x;
	input clk;
	input [31:0] A54x;
	input clk;
	input [31:0] A55x;
	input clk;
	input [31:0] A56x;
	input clk;
	input [31:0] A57x;
	input clk;
	input [31:0] A58x;
	input clk;
	input [31:0] A59x;
	input clk;
	input [31:0] A60x;
	input clk;
	input [31:0] A61x;
	input clk;
	input [31:0] A62x;
	input clk;
	input [31:0] A63x;
	input clk;
	input [31:0] A64x;
	input clk;
	input [31:0] A65x;
	input clk;
	input [31:0] A66x;
	input clk;
	input [31:0] A67x;
	input clk;
	input [31:0] A68x;
	input clk;
	input [31:0] A69x;
	input clk;
	input [31:0] A70x;
	input clk;
	input [31:0] A71x;
	input clk;
	input [31:0] A72x;
	input clk;
	input [31:0] A73x;
	input clk;
	input [31:0] A74x;
	input clk;
	input [31:0] A75x;
	input clk;
	input [31:0] A76x;
	input clk;
	input [31:0] A77x;
	input clk;
	input [31:0] A78x;
	input clk;
	input [31:0] A79x;
	input clk;
	input [31:0] A80x;
	input clk;
	input [31:0] A81x;
	input clk;
	input [31:0] A82x;
	input clk;
	input [31:0] A83x;
	input clk;
	input [31:0] A84x;
	input clk;
	input [31:0] A85x;
	input clk;
	input [31:0] A86x;
	input clk;
	input [31:0] A87x;
	input clk;
	input [31:0] A88x;
	input clk;
	input [31:0] A89x;
	input clk;
	input [31:0] A90x;
	input clk;
	input [31:0] A91x;
	input clk;
	input [31:0] A92x;
	input clk;
	input [31:0] A93x;
	input clk;
	input [31:0] A94x;
	input clk;
	input [31:0] A95x;
	input clk;
	input [31:0] A96x;
	input clk;
	input [31:0] A97x;
	input clk;
	input [31:0] A98x;
	input clk;
	input [31:0] A99x;
	input clk;
	input [31:0] A100x;
	input clk;
	input [31:0] A101x;
	input clk;
	input [31:0] A102x;
	input clk;
	input [31:0] A103x;
	input clk;
	input [31:0] A104x;
	input clk;
	input [31:0] A105x;
	input clk;
	input [31:0] A106x;
	input clk;
	input [31:0] A107x;
	input clk;
	input [31:0] A108x;
	input clk;
	input [31:0] A109x;
	input clk;
	input [31:0] A110x;
	input clk;
	input [31:0] A111x;
	input clk;
	input [31:0] A112x;
	input clk;
	input [31:0] A113x;
	input clk;
	input [31:0] A114x;
	input clk;
	input [31:0] A115x;
	input clk;
	input [31:0] A116x;
	input clk;
	input [31:0] A117x;
	input clk;
	input [31:0] A118x;
	input clk;
	input [31:0] A119x;
	input clk;
	input [31:0] A120x;
	input clk;
	input [31:0] A121x;
	input clk;
	input [31:0] A122x;
	input clk;
	input [31:0] A123x;
	input clk;
	input [31:0] A124x;
	input clk;
	input [31:0] A125x;
	input clk;
	input [31:0] A126x;
	input clk;
	input [31:0] A127x;
	input clk;
	input [31:0] A128x;
	input clk;
	input [31:0] A129x;
	input clk;
	input [31:0] A130x;
	input clk;
	input [31:0] A131x;
	input clk;
	input [31:0] A132x;
	input clk;
	input [31:0] A133x;
	input clk;
	input [31:0] A134x;
	input clk;
	input [31:0] A135x;
	input clk;
	input [31:0] A136x;
	input clk;
	input [31:0] A137x;
	input clk;
	input [31:0] A138x;
	input clk;
	input [31:0] A139x;
	input clk;
	input [31:0] A140x;
	input clk;
	input [31:0] A141x;
	input clk;
	input [31:0] A142x;
	input clk;
	input [31:0] A143x;
	input clk;
	input [31:0] A144x;
	input clk;
	input [31:0] A145x;
	input clk;
	input [31:0] A146x;
	input clk;
	input [31:0] A147x;
	input clk;
	input [31:0] A148x;
	input clk;
	input [31:0] A149x;
	input clk;
	input [31:0] A150x;
	input clk;
	input [31:0] A151x;
	input clk;
	input [31:0] A152x;
	input clk;
	input [31:0] A153x;
	input clk;
	input [31:0] A154x;
	input clk;
	input [31:0] A155x;
	input clk;
	input [31:0] A156x;
	input clk;
	input [31:0] A157x;
	input clk;
	input [31:0] A158x;
	input clk;
	input [31:0] A159x;
	input clk;
	input [31:0] A160x;
	input clk;
	input [31:0] A161x;
	input clk;
	input [31:0] A162x;
	input clk;
	input [31:0] A163x;
	input clk;
	input [31:0] A164x;
	input clk;
	input [31:0] A165x;
	input clk;
	input [31:0] A166x;
	input clk;
	input [31:0] A167x;
	input clk;
	input [31:0] A168x;
	input clk;
	input [31:0] A169x;
	input clk;
	input [31:0] A170x;
	input clk;
	input [31:0] A171x;
	input clk;
	input [31:0] A172x;
	input clk;
	input [31:0] A173x;
	input clk;
	input [31:0] A174x;
	input clk;
	input [31:0] A175x;
	input clk;
	input [31:0] A176x;
	input clk;
	input [31:0] A177x;
	input clk;
	input [31:0] A178x;
	input clk;
	input [31:0] A179x;
	input clk;
	input [31:0] A180x;
	input clk;
	input [31:0] A181x;
	input clk;
	input [31:0] A182x;
	input clk;
	input [31:0] A183x;
	input clk;
	input [31:0] A184x;
	input clk;
	input [31:0] A185x;
	input clk;
	input [31:0] A186x;
	output [31:0] N1x;
	reg [31:0] N1x; 

	parameter [31:0] W0x=32'b10111110010000100101111001110100;
	parameter [31:0] W1x=32'b00111110110010110100010001100101;
	parameter [31:0] W2x=32'b00111101010001011110101001100111;
	parameter [31:0] W3x=32'b10111110101111110111001100011011;
	parameter [31:0] W4x=32'b10111110001111011010010010100100;
	parameter [31:0] W5x=32'b10111101100111111101000100111101;
	parameter [31:0] W6x=32'b00111110110100111111101110000001;
	parameter [31:0] W7x=32'b00111101011010111100111010011000;
	parameter [31:0] W8x=32'b00111110110001111010110111100111;
	parameter [31:0] W9x=32'b00111110101010010011101110110010;
	parameter [31:0] W10x=32'b00111110100111100100010010110010;
	parameter [31:0] W11x=32'b00111110110000011111101000011000;
	parameter [31:0] W12x=32'b00111100111110000001010000100010;
	parameter [31:0] W13x=32'b10111011111001000101111000011000;
	parameter [31:0] W14x=32'b00111101111011100110000010110001;
	parameter [31:0] W15x=32'b10111100101000010110010010000010;
	parameter [31:0] W16x=32'b00111110000100000000110101011000;
	parameter [31:0] W17x=32'b10111110011001100011101010001010;
	parameter [31:0] W18x=32'b10111110001001000010100110011100;
	parameter [31:0] W19x=32'b00111100110011101101110011011100;
	parameter [31:0] W20x=32'b10111110001111000011011001101111;
	parameter [31:0] W21x=32'b00111110000001110110100111111000;
	parameter [31:0] W22x=32'b10111110001101111111110000000111;
	parameter [31:0] W23x=32'b10111101000010001001110110100000;
	parameter [31:0] W24x=32'b10111101100100000001001000011100;
	parameter [31:0] W25x=32'b10111110110011110101100010011111;
	parameter [31:0] W26x=32'b10111110110011111110010001110110;
	parameter [31:0] W27x=32'b10111110110111001000101101010101;
	parameter [31:0] W28x=32'b10111111000001100011011111000100;
	parameter [31:0] W29x=32'b10111110101110001001110000110011;
	parameter [31:0] W30x=32'b10111110100110110111010111001001;
	parameter [31:0] W31x=32'b10111110111011010011001000100111;
	parameter [31:0] W32x=32'b10111110011011101011001101001010;
	parameter [31:0] W33x=32'b10111110100100100000011001001111;
	parameter [31:0] W34x=32'b00111101001010000100100101100110;
	parameter [31:0] W35x=32'b00111011111101111001111001011000;
	parameter [31:0] W36x=32'b00111110011010110011011111010000;
	parameter [31:0] W37x=32'b10111100101100000011000111100010;
	parameter [31:0] W38x=32'b10111101100000110010110100101111;
	parameter [31:0] W39x=32'b10111100000010101010100111000011;
	parameter [31:0] W40x=32'b10111101001011000001110001010101;
	parameter [31:0] W41x=32'b00111101100010110101101101110000;
	parameter [31:0] W42x=32'b10111100110111101100001101100100;
	parameter [31:0] W43x=32'b00111101110011101010101010100100;
	parameter [31:0] W44x=32'b10111100010010010101101010101001;
	parameter [31:0] W45x=32'b10111100100101110000000111010001;
	parameter [31:0] W46x=32'b00111101110100010111111011101111;
	parameter [31:0] W47x=32'b00111101111111110110010000011011;
	parameter [31:0] W48x=32'b00111110100011011111001010000111;
	parameter [31:0] W49x=32'b00111110000110111101001100001000;
	parameter [31:0] W50x=32'b00111110001001110100001111110011;
	parameter [31:0] W51x=32'b00111101101000111110001011110100;
	parameter [31:0] W52x=32'b00111110001010111010101011011010;
	parameter [31:0] W53x=32'b00111101110111011010101001101100;
	parameter [31:0] W54x=32'b00111110010010011110101001011110;
	parameter [31:0] W55x=32'b00111101101100110001001101011011;
	parameter [31:0] W56x=32'b00111110010010100111111110110000;
	parameter [31:0] W57x=32'b00111110001010010011010111000111;
	parameter [31:0] W58x=32'b00111110100000100010100111110000;
	parameter [31:0] W59x=32'b00111110000110111010111010111010;
	parameter [31:0] W60x=32'b00111110100100001011100000100001;
	parameter [31:0] W61x=32'b00111110110010100010101000000100;
	parameter [31:0] W62x=32'b00111011000111001111001111110100;
	parameter [31:0] W63x=32'b00111110101101011011100010100111;
	parameter [31:0] W64x=32'b00111110000000101101001101001110;
	parameter [31:0] W65x=32'b00111110010001110100101000010110;
	parameter [31:0] W66x=32'b00111101111111011110000011000000;
	parameter [31:0] W67x=32'b00111110011010010101000110100010;
	parameter [31:0] W68x=32'b00111110001010101110011010100011;
	parameter [31:0] W69x=32'b00111101000110110100110001101101;
	parameter [31:0] W70x=32'b10111101110000001010110011001110;
	parameter [31:0] W71x=32'b00111101110111111101011111111001;
	parameter [31:0] W72x=32'b10111110010000110100011111111100;
	parameter [31:0] W73x=32'b10111110000001001111110001100110;
	parameter [31:0] W74x=32'b10111110000001100000011001001100;
	parameter [31:0] W75x=32'b10111110100001001000100001001000;
	parameter [31:0] W76x=32'b00111110000010110110110010100110;
	parameter [31:0] W77x=32'b00111011000000101001000011101001;
	parameter [31:0] W78x=32'b00111101101111001000001001100110;
	parameter [31:0] W79x=32'b00111101001011101110010010110110;
	parameter [31:0] W80x=32'b10111101000101110100111111010000;
	parameter [31:0] W81x=32'b00111110100111110110110001001010;
	parameter [31:0] W82x=32'b00111101000111010010001010100111;
	parameter [31:0] W83x=32'b00111110001101010110010010111001;
	parameter [31:0] W84x=32'b10111100111011010010000111011001;
	parameter [31:0] W85x=32'b10111110000001111100111001100110;
	parameter [31:0] W86x=32'b00111110101100010111100010000100;
	parameter [31:0] W87x=32'b10111110000011111000110001011111;
	parameter [31:0] W88x=32'b00111110000100101110110100110100;
	parameter [31:0] W89x=32'b00111100110100001110010001010000;
	parameter [31:0] W90x=32'b00111101111010011010101100110100;
	parameter [31:0] W91x=32'b00111101001100001101101111011010;
	parameter [31:0] W92x=32'b00111110000101011100111100100000;
	parameter [31:0] W93x=32'b00111101110100000010001100001111;
	parameter [31:0] W94x=32'b00111101111000000000010100110001;
	parameter [31:0] W95x=32'b00111101010110110101000100101111;
	parameter [31:0] W96x=32'b00111110011001001110101000001101;
	parameter [31:0] W97x=32'b10111101000000000010010100100111;
	parameter [31:0] W98x=32'b00111101110110011011000100000111;
	parameter [31:0] W99x=32'b00111101110001101111001010111100;
	parameter [31:0] W100x=32'b00111100011000001111000001110010;
	parameter [31:0] W101x=32'b00111101000001101101101110000110;
	parameter [31:0] W102x=32'b00111110001000010111000110011011;
	parameter [31:0] W103x=32'b00111110001101011100101001110010;
	parameter [31:0] W104x=32'b00111100001010000011100111101100;
	parameter [31:0] W105x=32'b00111101111111110101001100111110;
	parameter [31:0] W106x=32'b00111110100001100111110010110110;
	parameter [31:0] W107x=32'b10111110001001001100101011111100;
	parameter [31:0] W108x=32'b00111110010111001010011111101110;
	parameter [31:0] W109x=32'b00111101100110100101000001010101;
	parameter [31:0] W110x=32'b10111101100000100000100110110001;
	parameter [31:0] W111x=32'b00111101000000010111111101100110;
	parameter [31:0] W112x=32'b10111101100101110000011110100011;
	parameter [31:0] W113x=32'b00111110101001000110100001011010;
	parameter [31:0] W114x=32'b10111101001010100011000101110100;
	parameter [31:0] W115x=32'b10111101010111010110001000101001;
	parameter [31:0] W116x=32'b00111101110010111101000011011111;
	parameter [31:0] W117x=32'b00111101010110111111010000100100;
	parameter [31:0] W118x=32'b00111110001000010100011111011000;
	parameter [31:0] W119x=32'b00111011100110011101011110111110;
	parameter [31:0] W120x=32'b00111100101111110010010111101100;
	parameter [31:0] W121x=32'b00111110000011011001001101110111;
	parameter [31:0] W122x=32'b00111101100000101110000110011011;
	parameter [31:0] W123x=32'b00111101101110100100110100001110;
	parameter [31:0] W124x=32'b10111100011011010001001110001001;
	parameter [31:0] W125x=32'b00111101100110010110011010001110;
	parameter [31:0] W126x=32'b00111110001011110000000010010110;
	parameter [31:0] W127x=32'b10111101110110100101101010011110;
	parameter [31:0] W128x=32'b00111101101110111100111111010100;
	parameter [31:0] W129x=32'b00111101110111101001110001110111;
	parameter [31:0] W130x=32'b00111100011111101110110100110011;
	parameter [31:0] W131x=32'b00111110010010001000110011100000;
	parameter [31:0] W132x=32'b00111100110000100100001111000000;
	parameter [31:0] W133x=32'b00111101100001100100100001011111;
	parameter [31:0] W134x=32'b00111110000011000001011011010001;
	parameter [31:0] W135x=32'b10111101011001001000101101101001;
	parameter [31:0] W136x=32'b00111101111101101110000000101000;
	parameter [31:0] W137x=32'b00111110011000011100000001110001;
	parameter [31:0] W138x=32'b00111101110011110000110001110010;
	parameter [31:0] W139x=32'b10111101100101010001001100000101;
	parameter [31:0] W140x=32'b10111101011010000001101111110110;
	parameter [31:0] W141x=32'b00111110011000100101010100101100;
	parameter [31:0] W142x=32'b00111101010001000100000001110000;
	parameter [31:0] W143x=32'b10111110101100000001111011110100;
	parameter [31:0] W144x=32'b00111110010000010100000010111010;
	parameter [31:0] W145x=32'b10111101101110111000101111010101;
	parameter [31:0] W146x=32'b00111100011011010110000011101000;
	parameter [31:0] W147x=32'b00111110100111000111010110101111;
	parameter [31:0] W148x=32'b10111101111110100111000011100110;
	parameter [31:0] W149x=32'b00111110000001010000111110001001;
	parameter [31:0] W150x=32'b10111101001011110101110000111110;
	parameter [31:0] W151x=32'b00111101101101110011011100111110;
	parameter [31:0] W152x=32'b10111101101011110011111111110000;
	parameter [31:0] W153x=32'b00111110110101101001110000100010;
	parameter [31:0] W154x=32'b10111101010011111010111000001010;
	parameter [31:0] W155x=32'b00111101011110001100111000101100;
	parameter [31:0] W156x=32'b00111110010011010010100001000001;
	parameter [31:0] W157x=32'b00111101101100000110001000011100;
	parameter [31:0] W158x=32'b10111110100111001010010110000111;
	parameter [31:0] W159x=32'b10111100011110100001100110100001;
	parameter [31:0] W160x=32'b10111110000000010000001101110100;
	parameter [31:0] W161x=32'b00111110010111010111010010010010;
	parameter [31:0] W162x=32'b00111110001110000001001011000100;
	parameter [31:0] W163x=32'b10111110001110111111001000000010;
	parameter [31:0] W164x=32'b10111100101100110011001110000000;
	parameter [31:0] W165x=32'b00111110101100000101001110101101;
	parameter [31:0] W166x=32'b00111110101110000000001110110111;
	parameter [31:0] W167x=32'b10111101100001001011100010111001;
	parameter [31:0] W168x=32'b00111100111110100000101010010010;
	parameter [31:0] W169x=32'b00111110101100001000001000110100;
	parameter [31:0] W170x=32'b00111110100011100101011001100100;
	parameter [31:0] W171x=32'b00111110010100001110110101101000;
	parameter [31:0] W172x=32'b00111110111110100100101011101001;
	parameter [31:0] W173x=32'b10111101101010100001111100111001;
	parameter [31:0] W174x=32'b00111101100110100001000101110001;
	parameter [31:0] W175x=32'b10111101111011010111001101101110;
	parameter [31:0] W176x=32'b00111101101000100101110010011101;
	parameter [31:0] W177x=32'b10111110100001101101011010010111;
	parameter [31:0] W178x=32'b10111101010100100011001011100111;
	parameter [31:0] W179x=32'b00111101111101010010110110100110;
	parameter [31:0] W180x=32'b00111010000001111011001011111011;
	parameter [31:0] W181x=32'b00111110101000010001010100010000;
	parameter [31:0] W182x=32'b00111110101111010001111111010001;
	parameter [31:0] W183x=32'b10111111000001011011100000011010;
	parameter [31:0] W184x=32'b10111111000010011010011101101111;
	parameter [31:0] W185x=32'b10111111001111010000101110001001;
	parameter [31:0] W186x=32'b00111101100110111101000001011010;
	parameter [31:0] B0x=32'b10111100011110001100110010110000;
	wire [31:0] in0x;
	wire [31:0] in1x;
	wire [31:0] in2x;
	wire [31:0] in3x;
	wire [31:0] in4x;
	wire [31:0] in5x;
	wire [31:0] in6x;
	wire [31:0] in7x;
	wire [31:0] in8x;
	wire [31:0] in9x;
	wire [31:0] in10x;
	wire [31:0] in11x;
	wire [31:0] in12x;
	wire [31:0] in13x;
	wire [31:0] in14x;
	wire [31:0] in15x;
	wire [31:0] in16x;
	wire [31:0] in17x;
	wire [31:0] in18x;
	wire [31:0] in19x;
	wire [31:0] in20x;
	wire [31:0] in21x;
	wire [31:0] in22x;
	wire [31:0] in23x;
	wire [31:0] in24x;
	wire [31:0] in25x;
	wire [31:0] in26x;
	wire [31:0] in27x;
	wire [31:0] in28x;
	wire [31:0] in29x;
	wire [31:0] in30x;
	wire [31:0] in31x;
	wire [31:0] in32x;
	wire [31:0] in33x;
	wire [31:0] in34x;
	wire [31:0] in35x;
	wire [31:0] in36x;
	wire [31:0] in37x;
	wire [31:0] in38x;
	wire [31:0] in39x;
	wire [31:0] in40x;
	wire [31:0] in41x;
	wire [31:0] in42x;
	wire [31:0] in43x;
	wire [31:0] in44x;
	wire [31:0] in45x;
	wire [31:0] in46x;
	wire [31:0] in47x;
	wire [31:0] in48x;
	wire [31:0] in49x;
	wire [31:0] in50x;
	wire [31:0] in51x;
	wire [31:0] in52x;
	wire [31:0] in53x;
	wire [31:0] in54x;
	wire [31:0] in55x;
	wire [31:0] in56x;
	wire [31:0] in57x;
	wire [31:0] in58x;
	wire [31:0] in59x;
	wire [31:0] in60x;
	wire [31:0] in61x;
	wire [31:0] in62x;
	wire [31:0] in63x;
	wire [31:0] in64x;
	wire [31:0] in65x;
	wire [31:0] in66x;
	wire [31:0] in67x;
	wire [31:0] in68x;
	wire [31:0] in69x;
	wire [31:0] in70x;
	wire [31:0] in71x;
	wire [31:0] in72x;
	wire [31:0] in73x;
	wire [31:0] in74x;
	wire [31:0] in75x;
	wire [31:0] in76x;
	wire [31:0] in77x;
	wire [31:0] in78x;
	wire [31:0] in79x;
	wire [31:0] in80x;
	wire [31:0] in81x;
	wire [31:0] in82x;
	wire [31:0] in83x;
	wire [31:0] in84x;
	wire [31:0] in85x;
	wire [31:0] in86x;
	wire [31:0] in87x;
	wire [31:0] in88x;
	wire [31:0] in89x;
	wire [31:0] in90x;
	wire [31:0] in91x;
	wire [31:0] in92x;
	wire [31:0] in93x;
	wire [31:0] in94x;
	wire [31:0] in95x;
	wire [31:0] in96x;
	wire [31:0] in97x;
	wire [31:0] in98x;
	wire [31:0] in99x;
	wire [31:0] in100x;
	wire [31:0] in101x;
	wire [31:0] in102x;
	wire [31:0] in103x;
	wire [31:0] in104x;
	wire [31:0] in105x;
	wire [31:0] in106x;
	wire [31:0] in107x;
	wire [31:0] in108x;
	wire [31:0] in109x;
	wire [31:0] in110x;
	wire [31:0] in111x;
	wire [31:0] in112x;
	wire [31:0] in113x;
	wire [31:0] in114x;
	wire [31:0] in115x;
	wire [31:0] in116x;
	wire [31:0] in117x;
	wire [31:0] in118x;
	wire [31:0] in119x;
	wire [31:0] in120x;
	wire [31:0] in121x;
	wire [31:0] in122x;
	wire [31:0] in123x;
	wire [31:0] in124x;
	wire [31:0] in125x;
	wire [31:0] in126x;
	wire [31:0] in127x;
	wire [31:0] in128x;
	wire [31:0] in129x;
	wire [31:0] in130x;
	wire [31:0] in131x;
	wire [31:0] in132x;
	wire [31:0] in133x;
	wire [31:0] in134x;
	wire [31:0] in135x;
	wire [31:0] in136x;
	wire [31:0] in137x;
	wire [31:0] in138x;
	wire [31:0] in139x;
	wire [31:0] in140x;
	wire [31:0] in141x;
	wire [31:0] in142x;
	wire [31:0] in143x;
	wire [31:0] in144x;
	wire [31:0] in145x;
	wire [31:0] in146x;
	wire [31:0] in147x;
	wire [31:0] in148x;
	wire [31:0] in149x;
	wire [31:0] in150x;
	wire [31:0] in151x;
	wire [31:0] in152x;
	wire [31:0] in153x;
	wire [31:0] in154x;
	wire [31:0] in155x;
	wire [31:0] in156x;
	wire [31:0] in157x;
	wire [31:0] in158x;
	wire [31:0] in159x;
	wire [31:0] in160x;
	wire [31:0] in161x;
	wire [31:0] in162x;
	wire [31:0] in163x;
	wire [31:0] in164x;
	wire [31:0] in165x;
	wire [31:0] in166x;
	wire [31:0] in167x;
	wire [31:0] in168x;
	wire [31:0] in169x;
	wire [31:0] in170x;
	wire [31:0] in171x;
	wire [31:0] in172x;
	wire [31:0] in173x;
	wire [31:0] in174x;
	wire [31:0] in175x;
	wire [31:0] in176x;
	wire [31:0] in177x;
	wire [31:0] in178x;
	wire [31:0] in179x;
	wire [31:0] in180x;
	wire [31:0] in181x;
	wire [31:0] in182x;
	wire [31:0] in183x;
	wire [31:0] in184x;
	wire [31:0] in185x;
	wire [31:0] in186x;
	wire [31:0] sum0x;
	wire [31:0] sum1x;
	wire [31:0] sum2x;
	wire [31:0] sum3x;
	wire [31:0] sum4x;
	wire [31:0] sum5x;
	wire [31:0] sum6x;
	wire [31:0] sum7x;
	wire [31:0] sum8x;
	wire [31:0] sum9x;
	wire [31:0] sum10x;
	wire [31:0] sum11x;
	wire [31:0] sum12x;
	wire [31:0] sum13x;
	wire [31:0] sum14x;
	wire [31:0] sum15x;
	wire [31:0] sum16x;
	wire [31:0] sum17x;
	wire [31:0] sum18x;
	wire [31:0] sum19x;
	wire [31:0] sum20x;
	wire [31:0] sum21x;
	wire [31:0] sum22x;
	wire [31:0] sum23x;
	wire [31:0] sum24x;
	wire [31:0] sum25x;
	wire [31:0] sum26x;
	wire [31:0] sum27x;
	wire [31:0] sum28x;
	wire [31:0] sum29x;
	wire [31:0] sum30x;
	wire [31:0] sum31x;
	wire [31:0] sum32x;
	wire [31:0] sum33x;
	wire [31:0] sum34x;
	wire [31:0] sum35x;
	wire [31:0] sum36x;
	wire [31:0] sum37x;
	wire [31:0] sum38x;
	wire [31:0] sum39x;
	wire [31:0] sum40x;
	wire [31:0] sum41x;
	wire [31:0] sum42x;
	wire [31:0] sum43x;
	wire [31:0] sum44x;
	wire [31:0] sum45x;
	wire [31:0] sum46x;
	wire [31:0] sum47x;
	wire [31:0] sum48x;
	wire [31:0] sum49x;
	wire [31:0] sum50x;
	wire [31:0] sum51x;
	wire [31:0] sum52x;
	wire [31:0] sum53x;
	wire [31:0] sum54x;
	wire [31:0] sum55x;
	wire [31:0] sum56x;
	wire [31:0] sum57x;
	wire [31:0] sum58x;
	wire [31:0] sum59x;
	wire [31:0] sum60x;
	wire [31:0] sum61x;
	wire [31:0] sum62x;
	wire [31:0] sum63x;
	wire [31:0] sum64x;
	wire [31:0] sum65x;
	wire [31:0] sum66x;
	wire [31:0] sum67x;
	wire [31:0] sum68x;
	wire [31:0] sum69x;
	wire [31:0] sum70x;
	wire [31:0] sum71x;
	wire [31:0] sum72x;
	wire [31:0] sum73x;
	wire [31:0] sum74x;
	wire [31:0] sum75x;
	wire [31:0] sum76x;
	wire [31:0] sum77x;
	wire [31:0] sum78x;
	wire [31:0] sum79x;
	wire [31:0] sum80x;
	wire [31:0] sum81x;
	wire [31:0] sum82x;
	wire [31:0] sum83x;
	wire [31:0] sum84x;
	wire [31:0] sum85x;
	wire [31:0] sum86x;
	wire [31:0] sum87x;
	wire [31:0] sum88x;
	wire [31:0] sum89x;
	wire [31:0] sum90x;
	wire [31:0] sum91x;
	wire [31:0] sum92x;
	wire [31:0] sum93x;
	wire [31:0] sum94x;
	wire [31:0] sum95x;
	wire [31:0] sum96x;
	wire [31:0] sum97x;
	wire [31:0] sum98x;
	wire [31:0] sum99x;
	wire [31:0] sum100x;
	wire [31:0] sum101x;
	wire [31:0] sum102x;
	wire [31:0] sum103x;
	wire [31:0] sum104x;
	wire [31:0] sum105x;
	wire [31:0] sum106x;
	wire [31:0] sum107x;
	wire [31:0] sum108x;
	wire [31:0] sum109x;
	wire [31:0] sum110x;
	wire [31:0] sum111x;
	wire [31:0] sum112x;
	wire [31:0] sum113x;
	wire [31:0] sum114x;
	wire [31:0] sum115x;
	wire [31:0] sum116x;
	wire [31:0] sum117x;
	wire [31:0] sum118x;
	wire [31:0] sum119x;
	wire [31:0] sum120x;
	wire [31:0] sum121x;
	wire [31:0] sum122x;
	wire [31:0] sum123x;
	wire [31:0] sum124x;
	wire [31:0] sum125x;
	wire [31:0] sum126x;
	wire [31:0] sum127x;
	wire [31:0] sum128x;
	wire [31:0] sum129x;
	wire [31:0] sum130x;
	wire [31:0] sum131x;
	wire [31:0] sum132x;
	wire [31:0] sum133x;
	wire [31:0] sum134x;
	wire [31:0] sum135x;
	wire [31:0] sum136x;
	wire [31:0] sum137x;
	wire [31:0] sum138x;
	wire [31:0] sum139x;
	wire [31:0] sum140x;
	wire [31:0] sum141x;
	wire [31:0] sum142x;
	wire [31:0] sum143x;
	wire [31:0] sum144x;
	wire [31:0] sum145x;
	wire [31:0] sum146x;
	wire [31:0] sum147x;
	wire [31:0] sum148x;
	wire [31:0] sum149x;
	wire [31:0] sum150x;
	wire [31:0] sum151x;
	wire [31:0] sum152x;
	wire [31:0] sum153x;
	wire [31:0] sum154x;
	wire [31:0] sum155x;
	wire [31:0] sum156x;
	wire [31:0] sum157x;
	wire [31:0] sum158x;
	wire [31:0] sum159x;
	wire [31:0] sum160x;
	wire [31:0] sum161x;
	wire [31:0] sum162x;
	wire [31:0] sum163x;
	wire [31:0] sum164x;
	wire [31:0] sum165x;
	wire [31:0] sum166x;
	wire [31:0] sum167x;
	wire [31:0] sum168x;
	wire [31:0] sum169x;
	wire [31:0] sum170x;
	wire [31:0] sum171x;
	wire [31:0] sum172x;
	wire [31:0] sum173x;
	wire [31:0] sum174x;
	wire [31:0] sum175x;
	wire [31:0] sum176x;
	wire [31:0] sum177x;
	wire [31:0] sum178x;
	wire [31:0] sum179x;
	wire [31:0] sum180x;
	wire [31:0] sum181x;
	wire [31:0] sum182x;
	wire [31:0] sum183x;
	wire [31:0] sum184x;
	wire [31:0] sum185x;

	wire [31:0] sumout;
	float_mult mult0(
		.x(A0x),
		.y(W0x),
		.z(in0x));
	float_mult mult1(
		.x(A1x),
		.y(W1x),
		.z(in1x));
	float_mult mult2(
		.x(A2x),
		.y(W2x),
		.z(in2x));
	float_mult mult3(
		.x(A3x),
		.y(W3x),
		.z(in3x));
	float_mult mult4(
		.x(A4x),
		.y(W4x),
		.z(in4x));
	float_mult mult5(
		.x(A5x),
		.y(W5x),
		.z(in5x));
	float_mult mult6(
		.x(A6x),
		.y(W6x),
		.z(in6x));
	float_mult mult7(
		.x(A7x),
		.y(W7x),
		.z(in7x));
	float_mult mult8(
		.x(A8x),
		.y(W8x),
		.z(in8x));
	float_mult mult9(
		.x(A9x),
		.y(W9x),
		.z(in9x));
	float_mult mult10(
		.x(A10x),
		.y(W10x),
		.z(in10x));
	float_mult mult11(
		.x(A11x),
		.y(W11x),
		.z(in11x));
	float_mult mult12(
		.x(A12x),
		.y(W12x),
		.z(in12x));
	float_mult mult13(
		.x(A13x),
		.y(W13x),
		.z(in13x));
	float_mult mult14(
		.x(A14x),
		.y(W14x),
		.z(in14x));
	float_mult mult15(
		.x(A15x),
		.y(W15x),
		.z(in15x));
	float_mult mult16(
		.x(A16x),
		.y(W16x),
		.z(in16x));
	float_mult mult17(
		.x(A17x),
		.y(W17x),
		.z(in17x));
	float_mult mult18(
		.x(A18x),
		.y(W18x),
		.z(in18x));
	float_mult mult19(
		.x(A19x),
		.y(W19x),
		.z(in19x));
	float_mult mult20(
		.x(A20x),
		.y(W20x),
		.z(in20x));
	float_mult mult21(
		.x(A21x),
		.y(W21x),
		.z(in21x));
	float_mult mult22(
		.x(A22x),
		.y(W22x),
		.z(in22x));
	float_mult mult23(
		.x(A23x),
		.y(W23x),
		.z(in23x));
	float_mult mult24(
		.x(A24x),
		.y(W24x),
		.z(in24x));
	float_mult mult25(
		.x(A25x),
		.y(W25x),
		.z(in25x));
	float_mult mult26(
		.x(A26x),
		.y(W26x),
		.z(in26x));
	float_mult mult27(
		.x(A27x),
		.y(W27x),
		.z(in27x));
	float_mult mult28(
		.x(A28x),
		.y(W28x),
		.z(in28x));
	float_mult mult29(
		.x(A29x),
		.y(W29x),
		.z(in29x));
	float_mult mult30(
		.x(A30x),
		.y(W30x),
		.z(in30x));
	float_mult mult31(
		.x(A31x),
		.y(W31x),
		.z(in31x));
	float_mult mult32(
		.x(A32x),
		.y(W32x),
		.z(in32x));
	float_mult mult33(
		.x(A33x),
		.y(W33x),
		.z(in33x));
	float_mult mult34(
		.x(A34x),
		.y(W34x),
		.z(in34x));
	float_mult mult35(
		.x(A35x),
		.y(W35x),
		.z(in35x));
	float_mult mult36(
		.x(A36x),
		.y(W36x),
		.z(in36x));
	float_mult mult37(
		.x(A37x),
		.y(W37x),
		.z(in37x));
	float_mult mult38(
		.x(A38x),
		.y(W38x),
		.z(in38x));
	float_mult mult39(
		.x(A39x),
		.y(W39x),
		.z(in39x));
	float_mult mult40(
		.x(A40x),
		.y(W40x),
		.z(in40x));
	float_mult mult41(
		.x(A41x),
		.y(W41x),
		.z(in41x));
	float_mult mult42(
		.x(A42x),
		.y(W42x),
		.z(in42x));
	float_mult mult43(
		.x(A43x),
		.y(W43x),
		.z(in43x));
	float_mult mult44(
		.x(A44x),
		.y(W44x),
		.z(in44x));
	float_mult mult45(
		.x(A45x),
		.y(W45x),
		.z(in45x));
	float_mult mult46(
		.x(A46x),
		.y(W46x),
		.z(in46x));
	float_mult mult47(
		.x(A47x),
		.y(W47x),
		.z(in47x));
	float_mult mult48(
		.x(A48x),
		.y(W48x),
		.z(in48x));
	float_mult mult49(
		.x(A49x),
		.y(W49x),
		.z(in49x));
	float_mult mult50(
		.x(A50x),
		.y(W50x),
		.z(in50x));
	float_mult mult51(
		.x(A51x),
		.y(W51x),
		.z(in51x));
	float_mult mult52(
		.x(A52x),
		.y(W52x),
		.z(in52x));
	float_mult mult53(
		.x(A53x),
		.y(W53x),
		.z(in53x));
	float_mult mult54(
		.x(A54x),
		.y(W54x),
		.z(in54x));
	float_mult mult55(
		.x(A55x),
		.y(W55x),
		.z(in55x));
	float_mult mult56(
		.x(A56x),
		.y(W56x),
		.z(in56x));
	float_mult mult57(
		.x(A57x),
		.y(W57x),
		.z(in57x));
	float_mult mult58(
		.x(A58x),
		.y(W58x),
		.z(in58x));
	float_mult mult59(
		.x(A59x),
		.y(W59x),
		.z(in59x));
	float_mult mult60(
		.x(A60x),
		.y(W60x),
		.z(in60x));
	float_mult mult61(
		.x(A61x),
		.y(W61x),
		.z(in61x));
	float_mult mult62(
		.x(A62x),
		.y(W62x),
		.z(in62x));
	float_mult mult63(
		.x(A63x),
		.y(W63x),
		.z(in63x));
	float_mult mult64(
		.x(A64x),
		.y(W64x),
		.z(in64x));
	float_mult mult65(
		.x(A65x),
		.y(W65x),
		.z(in65x));
	float_mult mult66(
		.x(A66x),
		.y(W66x),
		.z(in66x));
	float_mult mult67(
		.x(A67x),
		.y(W67x),
		.z(in67x));
	float_mult mult68(
		.x(A68x),
		.y(W68x),
		.z(in68x));
	float_mult mult69(
		.x(A69x),
		.y(W69x),
		.z(in69x));
	float_mult mult70(
		.x(A70x),
		.y(W70x),
		.z(in70x));
	float_mult mult71(
		.x(A71x),
		.y(W71x),
		.z(in71x));
	float_mult mult72(
		.x(A72x),
		.y(W72x),
		.z(in72x));
	float_mult mult73(
		.x(A73x),
		.y(W73x),
		.z(in73x));
	float_mult mult74(
		.x(A74x),
		.y(W74x),
		.z(in74x));
	float_mult mult75(
		.x(A75x),
		.y(W75x),
		.z(in75x));
	float_mult mult76(
		.x(A76x),
		.y(W76x),
		.z(in76x));
	float_mult mult77(
		.x(A77x),
		.y(W77x),
		.z(in77x));
	float_mult mult78(
		.x(A78x),
		.y(W78x),
		.z(in78x));
	float_mult mult79(
		.x(A79x),
		.y(W79x),
		.z(in79x));
	float_mult mult80(
		.x(A80x),
		.y(W80x),
		.z(in80x));
	float_mult mult81(
		.x(A81x),
		.y(W81x),
		.z(in81x));
	float_mult mult82(
		.x(A82x),
		.y(W82x),
		.z(in82x));
	float_mult mult83(
		.x(A83x),
		.y(W83x),
		.z(in83x));
	float_mult mult84(
		.x(A84x),
		.y(W84x),
		.z(in84x));
	float_mult mult85(
		.x(A85x),
		.y(W85x),
		.z(in85x));
	float_mult mult86(
		.x(A86x),
		.y(W86x),
		.z(in86x));
	float_mult mult87(
		.x(A87x),
		.y(W87x),
		.z(in87x));
	float_mult mult88(
		.x(A88x),
		.y(W88x),
		.z(in88x));
	float_mult mult89(
		.x(A89x),
		.y(W89x),
		.z(in89x));
	float_mult mult90(
		.x(A90x),
		.y(W90x),
		.z(in90x));
	float_mult mult91(
		.x(A91x),
		.y(W91x),
		.z(in91x));
	float_mult mult92(
		.x(A92x),
		.y(W92x),
		.z(in92x));
	float_mult mult93(
		.x(A93x),
		.y(W93x),
		.z(in93x));
	float_mult mult94(
		.x(A94x),
		.y(W94x),
		.z(in94x));
	float_mult mult95(
		.x(A95x),
		.y(W95x),
		.z(in95x));
	float_mult mult96(
		.x(A96x),
		.y(W96x),
		.z(in96x));
	float_mult mult97(
		.x(A97x),
		.y(W97x),
		.z(in97x));
	float_mult mult98(
		.x(A98x),
		.y(W98x),
		.z(in98x));
	float_mult mult99(
		.x(A99x),
		.y(W99x),
		.z(in99x));
	float_mult mult100(
		.x(A100x),
		.y(W100x),
		.z(in100x));
	float_mult mult101(
		.x(A101x),
		.y(W101x),
		.z(in101x));
	float_mult mult102(
		.x(A102x),
		.y(W102x),
		.z(in102x));
	float_mult mult103(
		.x(A103x),
		.y(W103x),
		.z(in103x));
	float_mult mult104(
		.x(A104x),
		.y(W104x),
		.z(in104x));
	float_mult mult105(
		.x(A105x),
		.y(W105x),
		.z(in105x));
	float_mult mult106(
		.x(A106x),
		.y(W106x),
		.z(in106x));
	float_mult mult107(
		.x(A107x),
		.y(W107x),
		.z(in107x));
	float_mult mult108(
		.x(A108x),
		.y(W108x),
		.z(in108x));
	float_mult mult109(
		.x(A109x),
		.y(W109x),
		.z(in109x));
	float_mult mult110(
		.x(A110x),
		.y(W110x),
		.z(in110x));
	float_mult mult111(
		.x(A111x),
		.y(W111x),
		.z(in111x));
	float_mult mult112(
		.x(A112x),
		.y(W112x),
		.z(in112x));
	float_mult mult113(
		.x(A113x),
		.y(W113x),
		.z(in113x));
	float_mult mult114(
		.x(A114x),
		.y(W114x),
		.z(in114x));
	float_mult mult115(
		.x(A115x),
		.y(W115x),
		.z(in115x));
	float_mult mult116(
		.x(A116x),
		.y(W116x),
		.z(in116x));
	float_mult mult117(
		.x(A117x),
		.y(W117x),
		.z(in117x));
	float_mult mult118(
		.x(A118x),
		.y(W118x),
		.z(in118x));
	float_mult mult119(
		.x(A119x),
		.y(W119x),
		.z(in119x));
	float_mult mult120(
		.x(A120x),
		.y(W120x),
		.z(in120x));
	float_mult mult121(
		.x(A121x),
		.y(W121x),
		.z(in121x));
	float_mult mult122(
		.x(A122x),
		.y(W122x),
		.z(in122x));
	float_mult mult123(
		.x(A123x),
		.y(W123x),
		.z(in123x));
	float_mult mult124(
		.x(A124x),
		.y(W124x),
		.z(in124x));
	float_mult mult125(
		.x(A125x),
		.y(W125x),
		.z(in125x));
	float_mult mult126(
		.x(A126x),
		.y(W126x),
		.z(in126x));
	float_mult mult127(
		.x(A127x),
		.y(W127x),
		.z(in127x));
	float_mult mult128(
		.x(A128x),
		.y(W128x),
		.z(in128x));
	float_mult mult129(
		.x(A129x),
		.y(W129x),
		.z(in129x));
	float_mult mult130(
		.x(A130x),
		.y(W130x),
		.z(in130x));
	float_mult mult131(
		.x(A131x),
		.y(W131x),
		.z(in131x));
	float_mult mult132(
		.x(A132x),
		.y(W132x),
		.z(in132x));
	float_mult mult133(
		.x(A133x),
		.y(W133x),
		.z(in133x));
	float_mult mult134(
		.x(A134x),
		.y(W134x),
		.z(in134x));
	float_mult mult135(
		.x(A135x),
		.y(W135x),
		.z(in135x));
	float_mult mult136(
		.x(A136x),
		.y(W136x),
		.z(in136x));
	float_mult mult137(
		.x(A137x),
		.y(W137x),
		.z(in137x));
	float_mult mult138(
		.x(A138x),
		.y(W138x),
		.z(in138x));
	float_mult mult139(
		.x(A139x),
		.y(W139x),
		.z(in139x));
	float_mult mult140(
		.x(A140x),
		.y(W140x),
		.z(in140x));
	float_mult mult141(
		.x(A141x),
		.y(W141x),
		.z(in141x));
	float_mult mult142(
		.x(A142x),
		.y(W142x),
		.z(in142x));
	float_mult mult143(
		.x(A143x),
		.y(W143x),
		.z(in143x));
	float_mult mult144(
		.x(A144x),
		.y(W144x),
		.z(in144x));
	float_mult mult145(
		.x(A145x),
		.y(W145x),
		.z(in145x));
	float_mult mult146(
		.x(A146x),
		.y(W146x),
		.z(in146x));
	float_mult mult147(
		.x(A147x),
		.y(W147x),
		.z(in147x));
	float_mult mult148(
		.x(A148x),
		.y(W148x),
		.z(in148x));
	float_mult mult149(
		.x(A149x),
		.y(W149x),
		.z(in149x));
	float_mult mult150(
		.x(A150x),
		.y(W150x),
		.z(in150x));
	float_mult mult151(
		.x(A151x),
		.y(W151x),
		.z(in151x));
	float_mult mult152(
		.x(A152x),
		.y(W152x),
		.z(in152x));
	float_mult mult153(
		.x(A153x),
		.y(W153x),
		.z(in153x));
	float_mult mult154(
		.x(A154x),
		.y(W154x),
		.z(in154x));
	float_mult mult155(
		.x(A155x),
		.y(W155x),
		.z(in155x));
	float_mult mult156(
		.x(A156x),
		.y(W156x),
		.z(in156x));
	float_mult mult157(
		.x(A157x),
		.y(W157x),
		.z(in157x));
	float_mult mult158(
		.x(A158x),
		.y(W158x),
		.z(in158x));
	float_mult mult159(
		.x(A159x),
		.y(W159x),
		.z(in159x));
	float_mult mult160(
		.x(A160x),
		.y(W160x),
		.z(in160x));
	float_mult mult161(
		.x(A161x),
		.y(W161x),
		.z(in161x));
	float_mult mult162(
		.x(A162x),
		.y(W162x),
		.z(in162x));
	float_mult mult163(
		.x(A163x),
		.y(W163x),
		.z(in163x));
	float_mult mult164(
		.x(A164x),
		.y(W164x),
		.z(in164x));
	float_mult mult165(
		.x(A165x),
		.y(W165x),
		.z(in165x));
	float_mult mult166(
		.x(A166x),
		.y(W166x),
		.z(in166x));
	float_mult mult167(
		.x(A167x),
		.y(W167x),
		.z(in167x));
	float_mult mult168(
		.x(A168x),
		.y(W168x),
		.z(in168x));
	float_mult mult169(
		.x(A169x),
		.y(W169x),
		.z(in169x));
	float_mult mult170(
		.x(A170x),
		.y(W170x),
		.z(in170x));
	float_mult mult171(
		.x(A171x),
		.y(W171x),
		.z(in171x));
	float_mult mult172(
		.x(A172x),
		.y(W172x),
		.z(in172x));
	float_mult mult173(
		.x(A173x),
		.y(W173x),
		.z(in173x));
	float_mult mult174(
		.x(A174x),
		.y(W174x),
		.z(in174x));
	float_mult mult175(
		.x(A175x),
		.y(W175x),
		.z(in175x));
	float_mult mult176(
		.x(A176x),
		.y(W176x),
		.z(in176x));
	float_mult mult177(
		.x(A177x),
		.y(W177x),
		.z(in177x));
	float_mult mult178(
		.x(A178x),
		.y(W178x),
		.z(in178x));
	float_mult mult179(
		.x(A179x),
		.y(W179x),
		.z(in179x));
	float_mult mult180(
		.x(A180x),
		.y(W180x),
		.z(in180x));
	float_mult mult181(
		.x(A181x),
		.y(W181x),
		.z(in181x));
	float_mult mult182(
		.x(A182x),
		.y(W182x),
		.z(in182x));
	float_mult mult183(
		.x(A183x),
		.y(W183x),
		.z(in183x));
	float_mult mult184(
		.x(A184x),
		.y(W184x),
		.z(in184x));
	float_mult mult185(
		.x(A185x),
		.y(W185x),
		.z(in185x));
	float_mult mult186(
		.x(A186x),
		.y(W186x),
		.z(in186x));

	float_adder add0(
		.a(in0x),
		.b(in1x),
		.Out(sum0x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add1(
		.a(in2x),
		.b(in3x),
		.Out(sum1x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add2(
		.a(in4x),
		.b(in5x),
		.Out(sum2x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add3(
		.a(in6x),
		.b(in7x),
		.Out(sum3x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add4(
		.a(in8x),
		.b(in9x),
		.Out(sum4x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add5(
		.a(in10x),
		.b(in11x),
		.Out(sum5x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add6(
		.a(in12x),
		.b(in13x),
		.Out(sum6x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add7(
		.a(in14x),
		.b(in15x),
		.Out(sum7x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add8(
		.a(in16x),
		.b(in17x),
		.Out(sum8x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add9(
		.a(in18x),
		.b(in19x),
		.Out(sum9x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add10(
		.a(in20x),
		.b(in21x),
		.Out(sum10x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add11(
		.a(in22x),
		.b(in23x),
		.Out(sum11x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add12(
		.a(in24x),
		.b(in25x),
		.Out(sum12x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add13(
		.a(in26x),
		.b(in27x),
		.Out(sum13x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add14(
		.a(in28x),
		.b(in29x),
		.Out(sum14x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add15(
		.a(in30x),
		.b(in31x),
		.Out(sum15x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add16(
		.a(in32x),
		.b(in33x),
		.Out(sum16x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add17(
		.a(in34x),
		.b(in35x),
		.Out(sum17x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add18(
		.a(in36x),
		.b(in37x),
		.Out(sum18x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add19(
		.a(in38x),
		.b(in39x),
		.Out(sum19x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add20(
		.a(in40x),
		.b(in41x),
		.Out(sum20x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add21(
		.a(in42x),
		.b(in43x),
		.Out(sum21x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add22(
		.a(in44x),
		.b(in45x),
		.Out(sum22x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add23(
		.a(in46x),
		.b(in47x),
		.Out(sum23x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add24(
		.a(in48x),
		.b(in49x),
		.Out(sum24x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add25(
		.a(in50x),
		.b(in51x),
		.Out(sum25x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add26(
		.a(in52x),
		.b(in53x),
		.Out(sum26x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add27(
		.a(in54x),
		.b(in55x),
		.Out(sum27x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add28(
		.a(in56x),
		.b(in57x),
		.Out(sum28x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add29(
		.a(in58x),
		.b(in59x),
		.Out(sum29x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add30(
		.a(in60x),
		.b(in61x),
		.Out(sum30x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add31(
		.a(in62x),
		.b(in63x),
		.Out(sum31x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add32(
		.a(in64x),
		.b(in65x),
		.Out(sum32x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add33(
		.a(in66x),
		.b(in67x),
		.Out(sum33x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add34(
		.a(in68x),
		.b(in69x),
		.Out(sum34x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add35(
		.a(in70x),
		.b(in71x),
		.Out(sum35x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add36(
		.a(in72x),
		.b(in73x),
		.Out(sum36x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add37(
		.a(in74x),
		.b(in75x),
		.Out(sum37x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add38(
		.a(in76x),
		.b(in77x),
		.Out(sum38x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add39(
		.a(in78x),
		.b(in79x),
		.Out(sum39x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add40(
		.a(in80x),
		.b(in81x),
		.Out(sum40x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add41(
		.a(in82x),
		.b(in83x),
		.Out(sum41x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add42(
		.a(in84x),
		.b(in85x),
		.Out(sum42x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add43(
		.a(in86x),
		.b(in87x),
		.Out(sum43x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add44(
		.a(in88x),
		.b(in89x),
		.Out(sum44x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add45(
		.a(in90x),
		.b(in91x),
		.Out(sum45x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add46(
		.a(in92x),
		.b(in93x),
		.Out(sum46x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add47(
		.a(in94x),
		.b(in95x),
		.Out(sum47x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add48(
		.a(in96x),
		.b(in97x),
		.Out(sum48x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add49(
		.a(in98x),
		.b(in99x),
		.Out(sum49x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add50(
		.a(in100x),
		.b(in101x),
		.Out(sum50x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add51(
		.a(in102x),
		.b(in103x),
		.Out(sum51x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add52(
		.a(in104x),
		.b(in105x),
		.Out(sum52x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add53(
		.a(in106x),
		.b(in107x),
		.Out(sum53x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add54(
		.a(in108x),
		.b(in109x),
		.Out(sum54x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add55(
		.a(in110x),
		.b(in111x),
		.Out(sum55x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add56(
		.a(in112x),
		.b(in113x),
		.Out(sum56x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add57(
		.a(in114x),
		.b(in115x),
		.Out(sum57x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add58(
		.a(in116x),
		.b(in117x),
		.Out(sum58x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add59(
		.a(in118x),
		.b(in119x),
		.Out(sum59x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add60(
		.a(in120x),
		.b(in121x),
		.Out(sum60x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add61(
		.a(in122x),
		.b(in123x),
		.Out(sum61x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add62(
		.a(in124x),
		.b(in125x),
		.Out(sum62x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add63(
		.a(in126x),
		.b(in127x),
		.Out(sum63x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add64(
		.a(in128x),
		.b(in129x),
		.Out(sum64x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add65(
		.a(in130x),
		.b(in131x),
		.Out(sum65x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add66(
		.a(in132x),
		.b(in133x),
		.Out(sum66x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add67(
		.a(in134x),
		.b(in135x),
		.Out(sum67x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add68(
		.a(in136x),
		.b(in137x),
		.Out(sum68x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add69(
		.a(in138x),
		.b(in139x),
		.Out(sum69x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add70(
		.a(in140x),
		.b(in141x),
		.Out(sum70x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add71(
		.a(in142x),
		.b(in143x),
		.Out(sum71x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add72(
		.a(in144x),
		.b(in145x),
		.Out(sum72x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add73(
		.a(in146x),
		.b(in147x),
		.Out(sum73x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add74(
		.a(in148x),
		.b(in149x),
		.Out(sum74x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add75(
		.a(in150x),
		.b(in151x),
		.Out(sum75x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add76(
		.a(in152x),
		.b(in153x),
		.Out(sum76x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add77(
		.a(in154x),
		.b(in155x),
		.Out(sum77x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add78(
		.a(in156x),
		.b(in157x),
		.Out(sum78x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add79(
		.a(in158x),
		.b(in159x),
		.Out(sum79x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add80(
		.a(in160x),
		.b(in161x),
		.Out(sum80x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add81(
		.a(in162x),
		.b(in163x),
		.Out(sum81x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add82(
		.a(in164x),
		.b(in165x),
		.Out(sum82x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add83(
		.a(in166x),
		.b(in167x),
		.Out(sum83x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add84(
		.a(in168x),
		.b(in169x),
		.Out(sum84x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add85(
		.a(in170x),
		.b(in171x),
		.Out(sum85x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add86(
		.a(in172x),
		.b(in173x),
		.Out(sum86x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add87(
		.a(in174x),
		.b(in175x),
		.Out(sum87x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add88(
		.a(in176x),
		.b(in177x),
		.Out(sum88x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add89(
		.a(in178x),
		.b(in179x),
		.Out(sum89x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add90(
		.a(in180x),
		.b(in181x),
		.Out(sum90x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add91(
		.a(in182x),
		.b(in183x),
		.Out(sum91x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add92(
		.a(in184x),
		.b(in185x),
		.Out(sum92x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add93(
		.a(in186x),
		.b(B0x),
		.Out(sum93x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add94(
		.a(sum0x),
		.b(sum1x),
		.Out(sum94x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add95(
		.a(sum2x),
		.b(sum3x),
		.Out(sum95x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add96(
		.a(sum4x),
		.b(sum5x),
		.Out(sum96x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add97(
		.a(sum6x),
		.b(sum7x),
		.Out(sum97x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add98(
		.a(sum8x),
		.b(sum9x),
		.Out(sum98x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add99(
		.a(sum10x),
		.b(sum11x),
		.Out(sum99x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add100(
		.a(sum12x),
		.b(sum13x),
		.Out(sum100x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add101(
		.a(sum14x),
		.b(sum15x),
		.Out(sum101x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add102(
		.a(sum16x),
		.b(sum17x),
		.Out(sum102x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add103(
		.a(sum18x),
		.b(sum19x),
		.Out(sum103x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add104(
		.a(sum20x),
		.b(sum21x),
		.Out(sum104x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add105(
		.a(sum22x),
		.b(sum23x),
		.Out(sum105x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add106(
		.a(sum24x),
		.b(sum25x),
		.Out(sum106x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add107(
		.a(sum26x),
		.b(sum27x),
		.Out(sum107x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add108(
		.a(sum28x),
		.b(sum29x),
		.Out(sum108x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add109(
		.a(sum30x),
		.b(sum31x),
		.Out(sum109x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add110(
		.a(sum32x),
		.b(sum33x),
		.Out(sum110x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add111(
		.a(sum34x),
		.b(sum35x),
		.Out(sum111x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add112(
		.a(sum36x),
		.b(sum37x),
		.Out(sum112x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add113(
		.a(sum38x),
		.b(sum39x),
		.Out(sum113x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add114(
		.a(sum40x),
		.b(sum41x),
		.Out(sum114x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add115(
		.a(sum42x),
		.b(sum43x),
		.Out(sum115x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add116(
		.a(sum44x),
		.b(sum45x),
		.Out(sum116x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add117(
		.a(sum46x),
		.b(sum47x),
		.Out(sum117x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add118(
		.a(sum48x),
		.b(sum49x),
		.Out(sum118x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add119(
		.a(sum50x),
		.b(sum51x),
		.Out(sum119x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add120(
		.a(sum52x),
		.b(sum53x),
		.Out(sum120x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add121(
		.a(sum54x),
		.b(sum55x),
		.Out(sum121x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add122(
		.a(sum56x),
		.b(sum57x),
		.Out(sum122x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add123(
		.a(sum58x),
		.b(sum59x),
		.Out(sum123x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add124(
		.a(sum60x),
		.b(sum61x),
		.Out(sum124x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add125(
		.a(sum62x),
		.b(sum63x),
		.Out(sum125x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add126(
		.a(sum64x),
		.b(sum65x),
		.Out(sum126x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add127(
		.a(sum66x),
		.b(sum67x),
		.Out(sum127x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add128(
		.a(sum68x),
		.b(sum69x),
		.Out(sum128x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add129(
		.a(sum70x),
		.b(sum71x),
		.Out(sum129x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add130(
		.a(sum72x),
		.b(sum73x),
		.Out(sum130x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add131(
		.a(sum74x),
		.b(sum75x),
		.Out(sum131x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add132(
		.a(sum76x),
		.b(sum77x),
		.Out(sum132x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add133(
		.a(sum78x),
		.b(sum79x),
		.Out(sum133x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add134(
		.a(sum80x),
		.b(sum81x),
		.Out(sum134x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add135(
		.a(sum82x),
		.b(sum83x),
		.Out(sum135x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add136(
		.a(sum84x),
		.b(sum85x),
		.Out(sum136x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add137(
		.a(sum86x),
		.b(sum87x),
		.Out(sum137x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add138(
		.a(sum88x),
		.b(sum89x),
		.Out(sum138x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add139(
		.a(sum90x),
		.b(sum91x),
		.Out(sum139x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add140(
		.a(sum92x),
		.b(sum93x),
		.Out(sum140x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add141(
		.a(sum94x),
		.b(sum95x),
		.Out(sum141x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add142(
		.a(sum96x),
		.b(sum97x),
		.Out(sum142x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add143(
		.a(sum98x),
		.b(sum99x),
		.Out(sum143x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add144(
		.a(sum100x),
		.b(sum101x),
		.Out(sum144x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add145(
		.a(sum102x),
		.b(sum103x),
		.Out(sum145x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add146(
		.a(sum104x),
		.b(sum105x),
		.Out(sum146x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add147(
		.a(sum106x),
		.b(sum107x),
		.Out(sum147x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add148(
		.a(sum108x),
		.b(sum109x),
		.Out(sum148x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add149(
		.a(sum110x),
		.b(sum111x),
		.Out(sum149x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add150(
		.a(sum112x),
		.b(sum113x),
		.Out(sum150x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add151(
		.a(sum114x),
		.b(sum115x),
		.Out(sum151x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add152(
		.a(sum116x),
		.b(sum117x),
		.Out(sum152x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add153(
		.a(sum118x),
		.b(sum119x),
		.Out(sum153x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add154(
		.a(sum120x),
		.b(sum121x),
		.Out(sum154x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add155(
		.a(sum122x),
		.b(sum123x),
		.Out(sum155x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add156(
		.a(sum124x),
		.b(sum125x),
		.Out(sum156x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add157(
		.a(sum126x),
		.b(sum127x),
		.Out(sum157x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add158(
		.a(sum128x),
		.b(sum129x),
		.Out(sum158x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add159(
		.a(sum130x),
		.b(sum131x),
		.Out(sum159x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add160(
		.a(sum132x),
		.b(sum133x),
		.Out(sum160x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add161(
		.a(sum134x),
		.b(sum135x),
		.Out(sum161x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add162(
		.a(sum136x),
		.b(sum137x),
		.Out(sum162x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add163(
		.a(sum138x),
		.b(sum139x),
		.Out(sum163x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add164(
		.a(sum141x),
		.b(sum142x),
		.Out(sum164x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add165(
		.a(sum143x),
		.b(sum144x),
		.Out(sum165x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add166(
		.a(sum145x),
		.b(sum146x),
		.Out(sum166x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add167(
		.a(sum147x),
		.b(sum148x),
		.Out(sum167x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add168(
		.a(sum149x),
		.b(sum150x),
		.Out(sum168x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add169(
		.a(sum151x),
		.b(sum152x),
		.Out(sum169x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add170(
		.a(sum153x),
		.b(sum154x),
		.Out(sum170x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add171(
		.a(sum155x),
		.b(sum156x),
		.Out(sum171x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add172(
		.a(sum157x),
		.b(sum158x),
		.Out(sum172x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add173(
		.a(sum159x),
		.b(sum160x),
		.Out(sum173x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add174(
		.a(sum161x),
		.b(sum162x),
		.Out(sum174x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add175(
		.a(sum163x),
		.b(sum140x),
		.Out(sum175x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add176(
		.a(sum164x),
		.b(sum165x),
		.Out(sum176x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add177(
		.a(sum166x),
		.b(sum167x),
		.Out(sum177x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add178(
		.a(sum168x),
		.b(sum169x),
		.Out(sum178x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add179(
		.a(sum170x),
		.b(sum171x),
		.Out(sum179x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add180(
		.a(sum172x),
		.b(sum173x),
		.Out(sum180x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add181(
		.a(sum174x),
		.b(sum175x),
		.Out(sum181x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add182(
		.a(sum176x),
		.b(sum177x),
		.Out(sum182x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add183(
		.a(sum178x),
		.b(sum179x),
		.Out(sum183x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add184(
		.a(sum180x),
		.b(sum181x),
		.Out(sum184x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add185(
		.a(sum182x),
		.b(sum183x),
		.Out(sum185x),
		.Out_test(),
		.shift(),
		.c_out());

	float_adder add186(
		.a(sum185x),
		.b(sum184x),
		.Out(sumout),
		.Out_test(),
		.shift(),
		.c_out());
always@(posedge clk)
	begin 
		if(sumout[31]==0)
			N1x=sumout;
		else
			N1x=32'd0;
	end
endmodule
