module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = -4639;
	I1x = 6489;
	I2x = 5110;
	I3x = 6762;
	I4x = 7015;
	I5x = 473;
	I6x = 3970;
	I7x = 7624;
	I8x = 401;
	I9x = 6383;
	I10x = -5334;
	I11x = -7173;
	I12x = 5372;
	I13x = -5171;
	I14x = -463;
	I15x = -6842;
	I16x = -6573;
	I17x = -4224;
	I18x = -7250;
	I19x = 1974;
	I20x = -7124;
	I21x = 6596;
	I22x = 858;
	I23x = 1478;
	I24x = -3348;
	I25x = 4788;
	I26x = 1890;
	I27x = 6662;
	I28x = 1204;
	I29x = -2004;
	I30x = 4701;
	I31x = -1736;
	I32x = -3176;
	I33x = 3167;
	I34x = 4452;
	I35x = 4288;
	I36x = -5183;
	I37x = 742;
	I38x = 5130;
	I39x = -7811;
	I40x = 4378;
	I41x = -4067;
	I42x = -1357;
	I43x = 4005;
	I44x = 4122;
	I45x = 3806;
	I46x = 888;
	I47x = -6076;
	I48x = -6883;
	I49x = -5217;
	I50x = -2248;
	I51x = 116;
	I52x = 4898;
	I53x = -6379;
	I54x = -6779;
	I55x = -4624;
	I56x = -6015;
	I57x = 5174;
	I58x = -7961;
	I59x = -2444;
	I60x = -3210;
	I61x = -5887;
	I62x = -2314;
	I63x = -3316;
	I64x = -4038;
	I65x = -5016;
	I66x = 6853;
	I67x = -3180;
	I68x = -2514;
	I69x = -6206;
	I70x = 2891;
	I71x = 6885;
	I72x = 4578;
	I73x = 6851;
	I74x = 1449;
	I75x = 4141;
	I76x = 6381;
	I77x = 1259;
	I78x = 1220;
	I79x = 5456;
	I80x = -1264;
	I81x = -4144;
	I82x = -595;
	I83x = -3538;
	I84x = -2719;
	I85x = -3088;
	I86x = -8115;
	I87x = -5905;
	I88x = -4580;
	I89x = -2856;
	I90x = -4841;
	I91x = -4149;
	I92x = -6339;
	I93x = 3910;
	I94x = 1420;
	I95x = 5891;
	I96x = -2844;
	I97x = 7022;
	I98x = -3957;
	I99x = 6168;
	I100x = 2562;
	I101x = 2515;
	I102x = -3944;
	I103x = -882;
	I104x = 5156;
	I105x = -4168;
	I106x = 6420;
	I107x = 6869;
	I108x = 7782;
	I109x = -7294;
	I110x = -76;
	I111x = 6823;
	I112x = -3499;
	I113x = -1084;
	I114x = -7754;
	I115x = 7665;
	I116x = -108;
	I117x = 7727;
	I118x = 5443;
	I119x = -5383;
	I120x = 4020;
	I121x = -6070;
	I122x = -7166;
	I123x = 227;
	I124x = 1639;
	I125x = -2445;
	I126x = -3273;
	I127x = 2727;
	I128x = 7879;
	I129x = 6303;
	I130x = -2864;
	I131x = 1142;
	I132x = 5587;
	I133x = -4819;
	I134x = 7309;
	I135x = -8009;
	I136x = 2578;
	I137x = 2824;
	I138x = 6244;
	I139x = 455;
	I140x = -1850;
	I141x = 4037;
	I142x = 5135;
	I143x = -3298;
	I144x = 5109;
	I145x = 3115;
	I146x = -2775;
	I147x = -4902;
	I148x = 7021;
	I149x = -4852;
	I150x = 5785;
	I151x = 3234;
	I152x = 2105;
	I153x = -3660;
	I154x = 4631;
	I155x = -4313;
	I156x = -5724;
	I157x = 6973;
	I158x = -6692;
	I159x = -3177;
	I160x = -6475;
	I161x = 6947;
	I162x = -1206;
	I163x = -5792;
	I164x = -6414;
	I165x = -119;
	I166x = 5991;
	I167x = 6207;
	I168x = -5484;
	I169x = 6518;
	I170x = 888;
	I171x = 5885;
	I172x = 6149;
	I173x = 4624;
	I174x = 2955;
	I175x = -1069;
	I176x = 3588;
	I177x = -6926;
	I178x = -3301;
	I179x = 7611;
	I180x = -5300;
	I181x = 4207;
	I182x = 5098;
	I183x = 7096;
	I184x = 2267;
	I185x = 465;
	I186x = 867;
	end
endmodule
[0.         0.1623471  1.01006952 1.03976597 0.        ] 

 [0, 1329, 8274, 8517, 0] 

 ['0000000000000000', '0000010100110001', '0010000001010010', '0010000101000101', '0000000000000000']
