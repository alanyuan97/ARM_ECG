module layer_5(reset,clk,N1x,N2x,N3x,N4x,N5x,N6x,N7x,N8x,N9x,N10x,N11x,N12x,N13x,N14x,N15x,R0x,R1x,R2x,R3x,R4x,R5x,R6x,R7x,R8x,R9x,R10x,R11x,R12x,R13x,R14x,R15x,R16x,R17x,R18x,R19x,R20x,R21x,R22x,R23x,R24x,R25x,R26x,R27x,R28x,R29x);
	input reset, clk; 
	output [7:0] N1x,N2x,N3x,N4x,N5x,N6x,N7x,N8x,N9x,N10x,N11x,N12x,N13x,N14x,N15x;
	input [7:0] R0x,R1x,R2x,R3x,R4x,R5x,R6x,R7x,R8x,R9x,R10x,R11x,R12x,R13x,R14x,R15x,R16x,R17x,R18x,R19x,R20x,R21x,R22x,R23x,R24x,R25x,R26x,R27x,R28x,R29x;

	node_5_1 node_5_1( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N1x(N1x) 
	); 
	node_5_2 node_5_2( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N2x(N2x) 
	); 
	node_5_3 node_5_3( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N3x(N3x) 
	); 
	node_5_4 node_5_4( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N4x(N4x) 
	); 
	node_5_5 node_5_5( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N5x(N5x) 
	); 
	node_5_6 node_5_6( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N6x(N6x) 
	); 
	node_5_7 node_5_7( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N7x(N7x) 
	); 
	node_5_8 node_5_8( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N8x(N8x) 
	); 
	node_5_9 node_5_9( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N9x(N9x) 
	); 
	node_5_10 node_5_10( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N10x(N10x) 
	); 
	node_5_11 node_5_11( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N11x(N11x) 
	); 
	node_5_12 node_5_12( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N12x(N12x) 
	); 
	node_5_13 node_5_13( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N13x(N13x) 
	); 
	node_5_14 node_5_14( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N14x(N14x) 
	); 
	node_5_15 node_5_15( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.A15x(R15x), 
		.A16x(R16x), 
		.A17x(R17x), 
		.A18x(R18x), 
		.A19x(R19x), 
		.A20x(R20x), 
		.A21x(R21x), 
		.A22x(R22x), 
		.A23x(R23x), 
		.A24x(R24x), 
		.A25x(R25x), 
		.A26x(R26x), 
		.A27x(R27x), 
		.A28x(R28x), 
		.A29x(R29x), 
		.clk(clk), 
		.reset(reset), 
		.N15x(N15x) 
	); 
endmodule
