module rom_input(EN,data_add,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	input [9:0]data_add;
	output reg [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	always@(EN)
		begin
		case(data_add)
			9b'0b00000000:begin
				I0x <= 8175;
				I1x <= 4726;
				I2x <= 2908;
				I3x <= 1327;
				I4x <= 1310;
				I5x <= 1433;
				I6x <= 1449;
				I7x <= 1384;
				I8x <= 1425;
				I9x <= 1384;
				I10x <= 1368;
				I11x <= 1400;
				I12x <= 1400;
				I13x <= 1449;
				I14x <= 1425;
				I15x <= 1433;
				I16x <= 1507;
				I17x <= 1540;
				I18x <= 1638;
				I19x <= 1662;
				I20x <= 1712;
				I21x <= 1835;
				I22x <= 1916;
				I23x <= 2072;
				I24x <= 2154;
				I25x <= 2260;
				I26x <= 2424;
				I27x <= 2498;
				I28x <= 2629;
				I29x <= 2654;
				I30x <= 2703;
				I31x <= 2760;
				I32x <= 2670;
				I33x <= 2564;
				I34x <= 2285;
				I35x <= 2072;
				I36x <= 1908;
				I37x <= 1712;
				I38x <= 1638;
				I39x <= 1507;
				I40x <= 1441;
				I41x <= 1441;
				I42x <= 1409;
				I43x <= 1441;
				I44x <= 1392;
				I45x <= 1376;
				I46x <= 1400;
				I47x <= 1384;
				I48x <= 1449;
				I49x <= 1409;
				I50x <= 1400;
				I51x <= 1409;
				I52x <= 1400;
				I53x <= 1458;
				I54x <= 1409;
				I55x <= 1400;
				I56x <= 1425;
				I57x <= 1400;
				I58x <= 1449;
				I59x <= 1392;
				I60x <= 1359;
				I61x <= 1359;
				I62x <= 1343;
				I63x <= 1376;
				I64x <= 1318;
				I65x <= 1302;
				I66x <= 1327;
				I67x <= 1310;
				I68x <= 1359;
				I69x <= 1318;
				I70x <= 1335;
				I71x <= 1482;
				I72x <= 1548;
				I73x <= 1654;
				I74x <= 1581;
				I75x <= 1613;
				I76x <= 1720;
				I77x <= 1761;
				I78x <= 1785;
				I79x <= 1646;
				I80x <= 1409;
				I81x <= 1310;
				I82x <= 1236;
				I83x <= 1236;
				I84x <= 1146;
				I85x <= 1105;
				I86x <= 1130;
				I87x <= 1089;
				I88x <= 1146;
				I89x <= 1114;
				I90x <= 1097;
				I91x <= 1105;
				I92x <= 958;
				I93x <= 0;
				I94x <= 165;
				I95x <= 1974;
				I96x <= 5021;
				I97x <= 8192;
				I98x <= 5545;
				I99x <= 3457;
				I100x <= 1638;
				I101x <= 1204;
				I102x <= 1384;
				I103x <= 1474;
				I104x <= 1318;
				I105x <= 1318;
				I106x <= 1343;
				I107x <= 1335;
				I108x <= 1400;
				I109x <= 1384;
				I110x <= 1417;
				I111x <= 1482;
				I112x <= 1482;
				I113x <= 1548;
				I114x <= 1548;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000001:begin
				I0x <= 8192;
				I1x <= 3407;
				I2x <= 1957;
				I3x <= 478;
				I4x <= 667;
				I5x <= 1441;
				I6x <= 1916;
				I7x <= 1957;
				I8x <= 2048;
				I9x <= 1982;
				I10x <= 2015;
				I11x <= 2064;
				I12x <= 2023;
				I13x <= 2170;
				I14x <= 2228;
				I15x <= 2260;
				I16x <= 2277;
				I17x <= 2269;
				I18x <= 2416;
				I19x <= 2449;
				I20x <= 2441;
				I21x <= 2523;
				I22x <= 2670;
				I23x <= 2752;
				I24x <= 2801;
				I25x <= 2908;
				I26x <= 2949;
				I27x <= 3080;
				I28x <= 3104;
				I29x <= 3112;
				I30x <= 3260;
				I31x <= 3358;
				I32x <= 3399;
				I33x <= 3342;
				I34x <= 3162;
				I35x <= 2998;
				I36x <= 2490;
				I37x <= 2342;
				I38x <= 2228;
				I39x <= 1933;
				I40x <= 1785;
				I41x <= 1818;
				I42x <= 1843;
				I43x <= 1875;
				I44x <= 1843;
				I45x <= 1802;
				I46x <= 1916;
				I47x <= 1892;
				I48x <= 1859;
				I49x <= 1851;
				I50x <= 1933;
				I51x <= 1916;
				I52x <= 1875;
				I53x <= 1957;
				I54x <= 1925;
				I55x <= 1875;
				I56x <= 1818;
				I57x <= 1687;
				I58x <= 1695;
				I59x <= 1802;
				I60x <= 1679;
				I61x <= 1720;
				I62x <= 1728;
				I63x <= 1679;
				I64x <= 1818;
				I65x <= 1736;
				I66x <= 1695;
				I67x <= 1662;
				I68x <= 1703;
				I69x <= 1695;
				I70x <= 1900;
				I71x <= 2236;
				I72x <= 2498;
				I73x <= 2662;
				I74x <= 2883;
				I75x <= 3104;
				I76x <= 2686;
				I77x <= 2138;
				I78x <= 2170;
				I79x <= 1933;
				I80x <= 1564;
				I81x <= 1474;
				I82x <= 1474;
				I83x <= 1384;
				I84x <= 1286;
				I85x <= 1343;
				I86x <= 1302;
				I87x <= 1417;
				I88x <= 1499;
				I89x <= 1531;
				I90x <= 1482;
				I91x <= 1548;
				I92x <= 2031;
				I93x <= 2375;
				I94x <= 4046;
				I95x <= 8044;
				I96x <= 5218;
				I97x <= 1867;
				I98x <= 1089;
				I99x <= 0;
				I100x <= 791;
				I101x <= 1589;
				I102x <= 1892;
				I103x <= 1933;
				I104x <= 1998;
				I105x <= 2039;
				I106x <= 2080;
				I107x <= 1998;
				I108x <= 2154;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000010:begin
				I0x <= 8192;
				I1x <= 6881;
				I2x <= 3522;
				I3x <= 1441;
				I4x <= 0;
				I5x <= 412;
				I6x <= 966;
				I7x <= 901;
				I8x <= 909;
				I9x <= 909;
				I10x <= 909;
				I11x <= 958;
				I12x <= 950;
				I13x <= 958;
				I14x <= 1040;
				I15x <= 1146;
				I16x <= 1155;
				I17x <= 1122;
				I18x <= 1228;
				I19x <= 1302;
				I20x <= 1277;
				I21x <= 1384;
				I22x <= 1466;
				I23x <= 1540;
				I24x <= 1589;
				I25x <= 1654;
				I26x <= 1875;
				I27x <= 2056;
				I28x <= 2220;
				I29x <= 2465;
				I30x <= 2613;
				I31x <= 2826;
				I32x <= 2957;
				I33x <= 3055;
				I34x <= 3121;
				I35x <= 3088;
				I36x <= 2981;
				I37x <= 2768;
				I38x <= 2498;
				I39x <= 2211;
				I40x <= 1949;
				I41x <= 1630;
				I42x <= 1474;
				I43x <= 1376;
				I44x <= 1261;
				I45x <= 1146;
				I46x <= 1073;
				I47x <= 1056;
				I48x <= 1048;
				I49x <= 925;
				I50x <= 950;
				I51x <= 991;
				I52x <= 991;
				I53x <= 991;
				I54x <= 933;
				I55x <= 909;
				I56x <= 999;
				I57x <= 1007;
				I58x <= 1015;
				I59x <= 1007;
				I60x <= 1032;
				I61x <= 1024;
				I62x <= 1015;
				I63x <= 1024;
				I64x <= 1056;
				I65x <= 991;
				I66x <= 1015;
				I67x <= 1032;
				I68x <= 917;
				I69x <= 966;
				I70x <= 983;
				I71x <= 991;
				I72x <= 917;
				I73x <= 942;
				I74x <= 933;
				I75x <= 1015;
				I76x <= 974;
				I77x <= 909;
				I78x <= 933;
				I79x <= 925;
				I80x <= 942;
				I81x <= 909;
				I82x <= 933;
				I83x <= 917;
				I84x <= 909;
				I85x <= 827;
				I86x <= 860;
				I87x <= 909;
				I88x <= 835;
				I89x <= 884;
				I90x <= 868;
				I91x <= 835;
				I92x <= 835;
				I93x <= 851;
				I94x <= 860;
				I95x <= 835;
				I96x <= 851;
				I97x <= 909;
				I98x <= 818;
				I99x <= 876;
				I100x <= 868;
				I101x <= 901;
				I102x <= 892;
				I103x <= 876;
				I104x <= 901;
				I105x <= 958;
				I106x <= 933;
				I107x <= 991;
				I108x <= 1114;
				I109x <= 1245;
				I110x <= 1384;
				I111x <= 1556;
				I112x <= 1859;
				I113x <= 1941;
				I114x <= 1990;
				I115x <= 2072;
				I116x <= 1933;
				I117x <= 1785;
				I118x <= 1695;
				I119x <= 1368;
				I120x <= 1056;
				I121x <= 901;
				I122x <= 876;
				I123x <= 868;
				I124x <= 827;
				I125x <= 860;
				I126x <= 759;
				I127x <= 659;
				I128x <= 1294;
				I129x <= 4177;
				I130x <= 7733;
				I131x <= 7462;
				I132x <= 5480;
				I133x <= 3153;
				I134x <= 1179;
				I135x <= 308;
				I136x <= 688;
				I137x <= 1212;
				I138x <= 1187;
				I139x <= 1138;
				I140x <= 1236;
				I141x <= 1171;
				I142x <= 1286;
				I143x <= 1327;
				I144x <= 1310;
				I145x <= 1343;
				I146x <= 1351;
				I147x <= 1359;
				I148x <= 1482;
				I149x <= 1507;
				I150x <= 1613;
				I151x <= 1589;
				I152x <= 1712;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000011:begin
				I0x <= 7667;
				I1x <= 6447;
				I2x <= 3588;
				I3x <= 1622;
				I4x <= 50;
				I5x <= 0;
				I6x <= 424;
				I7x <= 694;
				I8x <= 670;
				I9x <= 697;
				I10x <= 717;
				I11x <= 738;
				I12x <= 774;
				I13x <= 792;
				I14x <= 810;
				I15x <= 843;
				I16x <= 942;
				I17x <= 991;
				I18x <= 1040;
				I19x <= 1056;
				I20x <= 1163;
				I21x <= 1245;
				I22x <= 1286;
				I23x <= 1351;
				I24x <= 1449;
				I25x <= 1548;
				I26x <= 1703;
				I27x <= 1867;
				I28x <= 2048;
				I29x <= 2220;
				I30x <= 2433;
				I31x <= 2637;
				I32x <= 2826;
				I33x <= 2957;
				I34x <= 3006;
				I35x <= 3014;
				I36x <= 2949;
				I37x <= 2744;
				I38x <= 2514;
				I39x <= 2228;
				I40x <= 1925;
				I41x <= 1703;
				I42x <= 1531;
				I43x <= 1368;
				I44x <= 1253;
				I45x <= 1155;
				I46x <= 1089;
				I47x <= 1056;
				I48x <= 1015;
				I49x <= 1015;
				I50x <= 999;
				I51x <= 958;
				I52x <= 958;
				I53x <= 950;
				I54x <= 991;
				I55x <= 1024;
				I56x <= 1024;
				I57x <= 1015;
				I58x <= 1048;
				I59x <= 1040;
				I60x <= 1073;
				I61x <= 1064;
				I62x <= 1040;
				I63x <= 1024;
				I64x <= 1040;
				I65x <= 1081;
				I66x <= 1056;
				I67x <= 1056;
				I68x <= 1040;
				I69x <= 999;
				I70x <= 991;
				I71x <= 966;
				I72x <= 974;
				I73x <= 983;
				I74x <= 966;
				I75x <= 958;
				I76x <= 950;
				I77x <= 933;
				I78x <= 950;
				I79x <= 933;
				I80x <= 966;
				I81x <= 1089;
				I82x <= 1269;
				I83x <= 1425;
				I84x <= 1662;
				I85x <= 1892;
				I86x <= 1990;
				I87x <= 2129;
				I88x <= 2195;
				I89x <= 1990;
				I90x <= 1802;
				I91x <= 1736;
				I92x <= 1515;
				I93x <= 1122;
				I94x <= 909;
				I95x <= 901;
				I96x <= 851;
				I97x <= 788;
				I98x <= 801;
				I99x <= 759;
				I100x <= 590;
				I101x <= 884;
				I102x <= 1703;
				I103x <= 4997;
				I104x <= 8192;
				I105x <= 7823;
				I106x <= 4939;
				I107x <= 2441;
				I108x <= 715;
				I109x <= 349;
				I110x <= 804;
				I111x <= 1105;
				I112x <= 1081;
				I113x <= 1105;
				I114x <= 1155;
				I115x <= 1163;
				I116x <= 1187;
				I117x <= 1212;
				I118x <= 1212;
				I119x <= 1302;
				I120x <= 1359;
				I121x <= 1400;
				I122x <= 1433;
				I123x <= 1499;
				I124x <= 1515;
				I125x <= 1613;
				I126x <= 1695;
				I127x <= 1753;
				I128x <= 1843;
				I129x <= 1966;
				I130x <= 2080;
				I131x <= 2252;
				I132x <= 2424;
				I133x <= 2654;
				I134x <= 2850;
				I135x <= 3055;
				I136x <= 3153;
				I137x <= 3284;
				I138x <= 3350;
				I139x <= 3350;
				I140x <= 3284;
				I141x <= 3129;
				I142x <= 2883;
				I143x <= 2605;
				I144x <= 2293;
				I145x <= 2088;
				I146x <= 1859;
				I147x <= 1687;
				I148x <= 1556;
				I149x <= 1441;
				I150x <= 1343;
				I151x <= 1318;
				I152x <= 1261;
				I153x <= 1245;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000100:begin
				I0x <= 7708;
				I1x <= 4603;
				I2x <= 2940;
				I3x <= 1802;
				I4x <= 1925;
				I5x <= 2023;
				I6x <= 2007;
				I7x <= 1957;
				I8x <= 1982;
				I9x <= 1990;
				I10x <= 2007;
				I11x <= 2023;
				I12x <= 2048;
				I13x <= 2088;
				I14x <= 2097;
				I15x <= 2146;
				I16x <= 2162;
				I17x <= 2211;
				I18x <= 2293;
				I19x <= 2334;
				I20x <= 2400;
				I21x <= 2473;
				I22x <= 2547;
				I23x <= 2686;
				I24x <= 2809;
				I25x <= 2924;
				I26x <= 3039;
				I27x <= 3145;
				I28x <= 3227;
				I29x <= 3268;
				I30x <= 3309;
				I31x <= 3301;
				I32x <= 3227;
				I33x <= 3022;
				I34x <= 2777;
				I35x <= 2547;
				I36x <= 2351;
				I37x <= 2187;
				I38x <= 2080;
				I39x <= 2031;
				I40x <= 1949;
				I41x <= 1933;
				I42x <= 1933;
				I43x <= 1941;
				I44x <= 1933;
				I45x <= 1908;
				I46x <= 1900;
				I47x <= 1900;
				I48x <= 1925;
				I49x <= 1925;
				I50x <= 1908;
				I51x <= 1900;
				I52x <= 1892;
				I53x <= 1875;
				I54x <= 1908;
				I55x <= 1900;
				I56x <= 1875;
				I57x <= 1892;
				I58x <= 1875;
				I59x <= 1875;
				I60x <= 1859;
				I61x <= 1884;
				I62x <= 1859;
				I63x <= 1859;
				I64x <= 1843;
				I65x <= 1859;
				I66x <= 1843;
				I67x <= 1818;
				I68x <= 1818;
				I69x <= 1810;
				I70x <= 1794;
				I71x <= 1777;
				I72x <= 1785;
				I73x <= 1777;
				I74x <= 1777;
				I75x <= 1761;
				I76x <= 1753;
				I77x <= 1744;
				I78x <= 1744;
				I79x <= 1785;
				I80x <= 1892;
				I81x <= 1990;
				I82x <= 2039;
				I83x <= 2039;
				I84x <= 2113;
				I85x <= 2203;
				I86x <= 2252;
				I87x <= 2146;
				I88x <= 2088;
				I89x <= 1826;
				I90x <= 1687;
				I91x <= 1630;
				I92x <= 1581;
				I93x <= 1531;
				I94x <= 1507;
				I95x <= 1490;
				I96x <= 1490;
				I97x <= 1499;
				I98x <= 1482;
				I99x <= 1474;
				I100x <= 1482;
				I101x <= 1466;
				I102x <= 1097;
				I103x <= 0;
				I104x <= 1007;
				I105x <= 3112;
				I106x <= 6094;
				I107x <= 8192;
				I108x <= 4907;
				I109x <= 3112;
				I110x <= 1540;
				I111x <= 1597;
				I112x <= 1744;
				I113x <= 1720;
				I114x <= 1687;
				I115x <= 1662;
				I116x <= 1687;
				I117x <= 1712;
				I118x <= 1695;
				I119x <= 1744;
				I120x <= 1769;
				I121x <= 1794;
				I122x <= 1810;
				I123x <= 1843;
				I124x <= 1867;
				I125x <= 1908;
				I126x <= 1982;
				I127x <= 2056;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000101:begin
				I0x <= 8192;
				I1x <= 7192;
				I2x <= 4161;
				I3x <= 1728;
				I4x <= 1277;
				I5x <= 1236;
				I6x <= 1310;
				I7x <= 1433;
				I8x <= 1400;
				I9x <= 1400;
				I10x <= 1531;
				I11x <= 1302;
				I12x <= 1359;
				I13x <= 1523;
				I14x <= 1376;
				I15x <= 1392;
				I16x <= 1466;
				I17x <= 1597;
				I18x <= 1818;
				I19x <= 1622;
				I20x <= 1925;
				I21x <= 1851;
				I22x <= 2211;
				I23x <= 2285;
				I24x <= 2359;
				I25x <= 2662;
				I26x <= 2875;
				I27x <= 3055;
				I28x <= 3301;
				I29x <= 3571;
				I30x <= 4005;
				I31x <= 3964;
				I32x <= 4038;
				I33x <= 4317;
				I34x <= 4218;
				I35x <= 4366;
				I36x <= 3907;
				I37x <= 3416;
				I38x <= 3047;
				I39x <= 2719;
				I40x <= 2383;
				I41x <= 2539;
				I42x <= 2023;
				I43x <= 1916;
				I44x <= 1818;
				I45x <= 1785;
				I46x <= 1638;
				I47x <= 1540;
				I48x <= 1753;
				I49x <= 1622;
				I50x <= 1638;
				I51x <= 1679;
				I52x <= 1622;
				I53x <= 1605;
				I54x <= 1622;
				I55x <= 1654;
				I56x <= 1802;
				I57x <= 1777;
				I58x <= 1703;
				I59x <= 1671;
				I60x <= 1613;
				I61x <= 1687;
				I62x <= 2105;
				I63x <= 1605;
				I64x <= 1564;
				I65x <= 1589;
				I66x <= 1540;
				I67x <= 1564;
				I68x <= 1794;
				I69x <= 1736;
				I70x <= 1392;
				I71x <= 1622;
				I72x <= 1376;
				I73x <= 1433;
				I74x <= 1835;
				I75x <= 1368;
				I76x <= 1417;
				I77x <= 1433;
				I78x <= 1556;
				I79x <= 1417;
				I80x <= 1220;
				I81x <= 1245;
				I82x <= 1343;
				I83x <= 1384;
				I84x <= 1417;
				I85x <= 1769;
				I86x <= 1843;
				I87x <= 2260;
				I88x <= 2031;
				I89x <= 2310;
				I90x <= 2531;
				I91x <= 2342;
				I92x <= 1916;
				I93x <= 2088;
				I94x <= 1671;
				I95x <= 1245;
				I96x <= 1130;
				I97x <= 1032;
				I98x <= 1032;
				I99x <= 925;
				I100x <= 933;
				I101x <= 901;
				I102x <= 991;
				I103x <= 1261;
				I104x <= 942;
				I105x <= 0;
				I106x <= 140;
				I107x <= 4218;
				I108x <= 7561;
				I109x <= 6545;
				I110x <= 3235;
				I111x <= 1196;
				I112x <= 655;
				I113x <= 868;
				I114x <= 1040;
				I115x <= 1155;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000110:begin
				I0x <= 8126;
				I1x <= 7741;
				I2x <= 1753;
				I3x <= 257;
				I4x <= 0;
				I5x <= 295;
				I6x <= 1032;
				I7x <= 1204;
				I8x <= 1212;
				I9x <= 1236;
				I10x <= 1228;
				I11x <= 1236;
				I12x <= 1269;
				I13x <= 1335;
				I14x <= 1327;
				I15x <= 1335;
				I16x <= 1359;
				I17x <= 1441;
				I18x <= 1474;
				I19x <= 1449;
				I20x <= 1474;
				I21x <= 1556;
				I22x <= 1662;
				I23x <= 1744;
				I24x <= 1802;
				I25x <= 1941;
				I26x <= 2023;
				I27x <= 2080;
				I28x <= 2195;
				I29x <= 2441;
				I30x <= 2670;
				I31x <= 2899;
				I32x <= 3186;
				I33x <= 3424;
				I34x <= 3653;
				I35x <= 3784;
				I36x <= 3932;
				I37x <= 4038;
				I38x <= 3956;
				I39x <= 3751;
				I40x <= 3342;
				I41x <= 2908;
				I42x <= 2441;
				I43x <= 2056;
				I44x <= 1695;
				I45x <= 1376;
				I46x <= 1212;
				I47x <= 991;
				I48x <= 950;
				I49x <= 876;
				I50x <= 876;
				I51x <= 876;
				I52x <= 819;
				I53x <= 876;
				I54x <= 909;
				I55x <= 999;
				I56x <= 1024;
				I57x <= 1040;
				I58x <= 1015;
				I59x <= 1015;
				I60x <= 1015;
				I61x <= 1040;
				I62x <= 1081;
				I63x <= 1064;
				I64x <= 1081;
				I65x <= 1024;
				I66x <= 999;
				I67x <= 983;
				I68x <= 942;
				I69x <= 884;
				I70x <= 884;
				I71x <= 843;
				I72x <= 819;
				I73x <= 795;
				I74x <= 753;
				I75x <= 753;
				I76x <= 719;
				I77x <= 730;
				I78x <= 761;
				I79x <= 699;
				I80x <= 638;
				I81x <= 656;
				I82x <= 642;
				I83x <= 649;
				I84x <= 638;
				I85x <= 626;
				I86x <= 688;
				I87x <= 719;
				I88x <= 738;
				I89x <= 780;
				I90x <= 819;
				I91x <= 827;
				I92x <= 827;
				I93x <= 772;
				I94x <= 780;
				I95x <= 795;
				I96x <= 835;
				I97x <= 819;
				I98x <= 835;
				I99x <= 819;
				I100x <= 792;
				I101x <= 819;
				I102x <= 860;
				I103x <= 925;
				I104x <= 1204;
				I105x <= 1294;
				I106x <= 1458;
				I107x <= 1540;
				I108x <= 1671;
				I109x <= 1654;
				I110x <= 1572;
				I111x <= 1253;
				I112x <= 1204;
				I113x <= 1081;
				I114x <= 884;
				I115x <= 792;
				I116x <= 811;
				I117x <= 788;
				I118x <= 788;
				I119x <= 811;
				I120x <= 788;
				I121x <= 806;
				I122x <= 884;
				I123x <= 795;
				I124x <= 195;
				I125x <= 480;
				I126x <= 3563;
				I127x <= 7716;
				I128x <= 8192;
				I129x <= 2228;
				I130x <= 231;
				I131x <= 7;
				I132x <= 115;
				I133x <= 1015;
				I134x <= 1261;
				I135x <= 1269;
				I136x <= 1318;
				I137x <= 1318;
				I138x <= 1310;
				I139x <= 1351;
				I140x <= 1335;
				I141x <= 1466;
				I142x <= 1507;
				I143x <= 1523;
				I144x <= 1490;
				I145x <= 1540;
				I146x <= 1605;
				I147x <= 1671;
				I148x <= 1744;
				I149x <= 1761;
				I150x <= 1867;
				I151x <= 1892;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00000111:begin
				I0x <= 7954;
				I1x <= 6291;
				I2x <= 1703;
				I3x <= 0;
				I4x <= 217;
				I5x <= 1269;
				I6x <= 1802;
				I7x <= 1982;
				I8x <= 2072;
				I9x <= 2129;
				I10x <= 2154;
				I11x <= 2228;
				I12x <= 2269;
				I13x <= 2318;
				I14x <= 2318;
				I15x <= 2326;
				I16x <= 2342;
				I17x <= 2408;
				I18x <= 2457;
				I19x <= 2547;
				I20x <= 2564;
				I21x <= 2719;
				I22x <= 2867;
				I23x <= 2990;
				I24x <= 3121;
				I25x <= 3252;
				I26x <= 3416;
				I27x <= 3620;
				I28x <= 3883;
				I29x <= 4128;
				I30x <= 4382;
				I31x <= 4595;
				I32x <= 4775;
				I33x <= 4833;
				I34x <= 4734;
				I35x <= 4489;
				I36x <= 4112;
				I37x <= 3751;
				I38x <= 3399;
				I39x <= 3039;
				I40x <= 2744;
				I41x <= 2588;
				I42x <= 2473;
				I43x <= 2359;
				I44x <= 2375;
				I45x <= 2334;
				I46x <= 2293;
				I47x <= 2285;
				I48x <= 2203;
				I49x <= 2146;
				I50x <= 2113;
				I51x <= 2097;
				I52x <= 2113;
				I53x <= 2080;
				I54x <= 2097;
				I55x <= 2080;
				I56x <= 2138;
				I57x <= 2105;
				I58x <= 2121;
				I59x <= 2138;
				I60x <= 2146;
				I61x <= 2097;
				I62x <= 2080;
				I63x <= 2064;
				I64x <= 2064;
				I65x <= 2039;
				I66x <= 2048;
				I67x <= 2056;
				I68x <= 2072;
				I69x <= 2072;
				I70x <= 2105;
				I71x <= 2072;
				I72x <= 2048;
				I73x <= 2056;
				I74x <= 2121;
				I75x <= 2129;
				I76x <= 2080;
				I77x <= 2088;
				I78x <= 2056;
				I79x <= 2023;
				I80x <= 2015;
				I81x <= 1966;
				I82x <= 1949;
				I83x <= 1900;
				I84x <= 1933;
				I85x <= 1998;
				I86x <= 1974;
				I87x <= 1990;
				I88x <= 1998;
				I89x <= 1998;
				I90x <= 1957;
				I91x <= 1974;
				I92x <= 2015;
				I93x <= 2048;
				I94x <= 2056;
				I95x <= 2015;
				I96x <= 2056;
				I97x <= 2080;
				I98x <= 2072;
				I99x <= 2056;
				I100x <= 2023;
				I101x <= 1974;
				I102x <= 2064;
				I103x <= 2039;
				I104x <= 2023;
				I105x <= 2228;
				I106x <= 2473;
				I107x <= 2367;
				I108x <= 2367;
				I109x <= 2072;
				I110x <= 2146;
				I111x <= 2048;
				I112x <= 2064;
				I113x <= 1974;
				I114x <= 1957;
				I115x <= 1957;
				I116x <= 2056;
				I117x <= 2015;
				I118x <= 2056;
				I119x <= 2023;
				I120x <= 1974;
				I121x <= 1908;
				I122x <= 1744;
				I123x <= 2441;
				I124x <= 3850;
				I125x <= 5840;
				I126x <= 8192;
				I127x <= 6217;
				I128x <= 1925;
				I129x <= 402;
				I130x <= 729;
				I131x <= 1703;
				I132x <= 2154;
				I133x <= 2334;
				I134x <= 2351;
				I135x <= 2375;
				I136x <= 2441;
				I137x <= 2506;
				I138x <= 2506;
				I139x <= 2605;
				I140x <= 2646;
				I141x <= 2678;
				I142x <= 2670;
				I143x <= 2686;
				I144x <= 2711;
				I145x <= 2801;
				I146x <= 2875;
				I147x <= 2924;
				I148x <= 3006;
				I149x <= 3096;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001000:begin
				I0x <= 8019;
				I1x <= 7626;
				I2x <= 3956;
				I3x <= 0;
				I4x <= 1105;
				I5x <= 2260;
				I6x <= 3637;
				I7x <= 3063;
				I8x <= 2473;
				I9x <= 2744;
				I10x <= 2793;
				I11x <= 2662;
				I12x <= 2990;
				I13x <= 2859;
				I14x <= 3014;
				I15x <= 3178;
				I16x <= 3203;
				I17x <= 3383;
				I18x <= 3375;
				I19x <= 3497;
				I20x <= 3776;
				I21x <= 3833;
				I22x <= 4358;
				I23x <= 4407;
				I24x <= 5087;
				I25x <= 5054;
				I26x <= 5152;
				I27x <= 5603;
				I28x <= 5701;
				I29x <= 5668;
				I30x <= 5660;
				I31x <= 5611;
				I32x <= 5611;
				I33x <= 5177;
				I34x <= 4947;
				I35x <= 4300;
				I36x <= 4161;
				I37x <= 3866;
				I38x <= 3440;
				I39x <= 3629;
				I40x <= 3252;
				I41x <= 3129;
				I42x <= 3186;
				I43x <= 3121;
				I44x <= 3309;
				I45x <= 3145;
				I46x <= 3104;
				I47x <= 3252;
				I48x <= 3153;
				I49x <= 3276;
				I50x <= 3153;
				I51x <= 3219;
				I52x <= 3252;
				I53x <= 3219;
				I54x <= 3252;
				I55x <= 3211;
				I56x <= 3104;
				I57x <= 3801;
				I58x <= 3981;
				I59x <= 4210;
				I60x <= 4407;
				I61x <= 4620;
				I62x <= 4726;
				I63x <= 4751;
				I64x <= 4718;
				I65x <= 5062;
				I66x <= 4448;
				I67x <= 4186;
				I68x <= 3538;
				I69x <= 3211;
				I70x <= 2891;
				I71x <= 2727;
				I72x <= 2760;
				I73x <= 2572;
				I74x <= 2629;
				I75x <= 2433;
				I76x <= 2441;
				I77x <= 3047;
				I78x <= 3604;
				I79x <= 5873;
				I80x <= 8192;
				I81x <= 5521;
				I82x <= 1572;
				I83x <= 524;
				I84x <= 1277;
				I85x <= 3538;
				I86x <= 3088;
				I87x <= 2711;
				I88x <= 2695;
				I89x <= 2867;
				I90x <= 2744;
				I91x <= 2752;
				I92x <= 2908;
				I93x <= 2990;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001001:begin
				I0x <= 7774;
				I1x <= 7184;
				I2x <= 3948;
				I3x <= 1712;
				I4x <= 364;
				I5x <= 1736;
				I6x <= 2670;
				I7x <= 2809;
				I8x <= 2924;
				I9x <= 3014;
				I10x <= 3129;
				I11x <= 3211;
				I12x <= 3252;
				I13x <= 3268;
				I14x <= 3260;
				I15x <= 3203;
				I16x <= 3301;
				I17x <= 3432;
				I18x <= 3481;
				I19x <= 3538;
				I20x <= 3825;
				I21x <= 3760;
				I22x <= 3956;
				I23x <= 4235;
				I24x <= 4521;
				I25x <= 4808;
				I26x <= 5136;
				I27x <= 5505;
				I28x <= 5816;
				I29x <= 6094;
				I30x <= 6250;
				I31x <= 6381;
				I32x <= 6250;
				I33x <= 5881;
				I34x <= 5365;
				I35x <= 4767;
				I36x <= 4177;
				I37x <= 3653;
				I38x <= 3268;
				I39x <= 2891;
				I40x <= 2826;
				I41x <= 2736;
				I42x <= 2662;
				I43x <= 2588;
				I44x <= 2555;
				I45x <= 2605;
				I46x <= 2588;
				I47x <= 2498;
				I48x <= 2490;
				I49x <= 2531;
				I50x <= 2514;
				I51x <= 2547;
				I52x <= 2506;
				I53x <= 2572;
				I54x <= 2605;
				I55x <= 2621;
				I56x <= 2646;
				I57x <= 2629;
				I58x <= 2703;
				I59x <= 2678;
				I60x <= 2686;
				I61x <= 2686;
				I62x <= 2621;
				I63x <= 2588;
				I64x <= 2596;
				I65x <= 2588;
				I66x <= 2555;
				I67x <= 2588;
				I68x <= 2498;
				I69x <= 2564;
				I70x <= 2416;
				I71x <= 2449;
				I72x <= 2301;
				I73x <= 2342;
				I74x <= 2318;
				I75x <= 2260;
				I76x <= 2269;
				I77x <= 2228;
				I78x <= 2236;
				I79x <= 2277;
				I80x <= 2277;
				I81x <= 2244;
				I82x <= 2269;
				I83x <= 2228;
				I84x <= 2277;
				I85x <= 2260;
				I86x <= 2228;
				I87x <= 2220;
				I88x <= 2195;
				I89x <= 2260;
				I90x <= 2670;
				I91x <= 2891;
				I92x <= 2965;
				I93x <= 3276;
				I94x <= 3432;
				I95x <= 3055;
				I96x <= 3186;
				I97x <= 3284;
				I98x <= 2580;
				I99x <= 2416;
				I100x <= 2056;
				I101x <= 2048;
				I102x <= 2129;
				I103x <= 2064;
				I104x <= 2031;
				I105x <= 2007;
				I106x <= 2113;
				I107x <= 2039;
				I108x <= 2080;
				I109x <= 2875;
				I110x <= 3383;
				I111x <= 4079;
				I112x <= 7315;
				I113x <= 8192;
				I114x <= 5251;
				I115x <= 1974;
				I116x <= 0;
				I117x <= 892;
				I118x <= 2162;
				I119x <= 2416;
				I120x <= 2465;
				I121x <= 2654;
				I122x <= 2768;
				I123x <= 2859;
				I124x <= 2891;
				I125x <= 2973;
				I126x <= 3031;
				I127x <= 3006;
				I128x <= 3031;
				I129x <= 3096;
				I130x <= 3235;
				I131x <= 3293;
				I132x <= 3448;
				I133x <= 3571;
				I134x <= 3751;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001010:begin
				I0x <= 8192;
				I1x <= 6766;
				I2x <= 1925;
				I3x <= 152;
				I4x <= 473;
				I5x <= 1130;
				I6x <= 1015;
				I7x <= 958;
				I8x <= 925;
				I9x <= 884;
				I10x <= 892;
				I11x <= 917;
				I12x <= 925;
				I13x <= 966;
				I14x <= 983;
				I15x <= 966;
				I16x <= 983;
				I17x <= 958;
				I18x <= 991;
				I19x <= 1097;
				I20x <= 1130;
				I21x <= 1155;
				I22x <= 1236;
				I23x <= 1286;
				I24x <= 1376;
				I25x <= 1433;
				I26x <= 1556;
				I27x <= 1662;
				I28x <= 1843;
				I29x <= 2113;
				I30x <= 2334;
				I31x <= 2662;
				I32x <= 2883;
				I33x <= 3080;
				I34x <= 3301;
				I35x <= 3563;
				I36x <= 3588;
				I37x <= 3424;
				I38x <= 3022;
				I39x <= 2506;
				I40x <= 2048;
				I41x <= 1556;
				I42x <= 1269;
				I43x <= 1015;
				I44x <= 876;
				I45x <= 757;
				I46x <= 648;
				I47x <= 691;
				I48x <= 681;
				I49x <= 668;
				I50x <= 691;
				I51x <= 720;
				I52x <= 747;
				I53x <= 734;
				I54x <= 774;
				I55x <= 738;
				I56x <= 714;
				I57x <= 724;
				I58x <= 728;
				I59x <= 741;
				I60x <= 754;
				I61x <= 747;
				I62x <= 757;
				I63x <= 764;
				I64x <= 728;
				I65x <= 741;
				I66x <= 744;
				I67x <= 764;
				I68x <= 694;
				I69x <= 648;
				I70x <= 720;
				I71x <= 751;
				I72x <= 757;
				I73x <= 738;
				I74x <= 751;
				I75x <= 761;
				I76x <= 744;
				I77x <= 767;
				I78x <= 757;
				I79x <= 714;
				I80x <= 901;
				I81x <= 1064;
				I82x <= 1105;
				I83x <= 1073;
				I84x <= 1196;
				I85x <= 1212;
				I86x <= 1130;
				I87x <= 1064;
				I88x <= 925;
				I89x <= 884;
				I90x <= 764;
				I91x <= 655;
				I92x <= 595;
				I93x <= 535;
				I94x <= 535;
				I95x <= 506;
				I96x <= 502;
				I97x <= 529;
				I98x <= 522;
				I99x <= 562;
				I100x <= 545;
				I101x <= 512;
				I102x <= 449;
				I103x <= 0;
				I104x <= 158;
				I105x <= 1548;
				I106x <= 4997;
				I107x <= 7979;
				I108x <= 6356;
				I109x <= 1687;
				I110x <= 165;
				I111x <= 443;
				I112x <= 1015;
				I113x <= 950;
				I114x <= 843;
				I115x <= 800;
				I116x <= 827;
				I117x <= 827;
				I118x <= 843;
				I119x <= 851;
				I120x <= 827;
				I121x <= 843;
				I122x <= 827;
				I123x <= 892;
				I124x <= 892;
				I125x <= 925;
				I126x <= 958;
				I127x <= 1032;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001011:begin
				I0x <= 7897;
				I1x <= 3874;
				I2x <= 1916;
				I3x <= 185;
				I4x <= 0;
				I5x <= 725;
				I6x <= 1261;
				I7x <= 1482;
				I8x <= 1425;
				I9x <= 1556;
				I10x <= 1564;
				I11x <= 1662;
				I12x <= 1622;
				I13x <= 1671;
				I14x <= 1638;
				I15x <= 1712;
				I16x <= 1753;
				I17x <= 1851;
				I18x <= 1867;
				I19x <= 1908;
				I20x <= 2064;
				I21x <= 2097;
				I22x <= 2310;
				I23x <= 2359;
				I24x <= 2506;
				I25x <= 2629;
				I26x <= 2736;
				I27x <= 2867;
				I28x <= 2940;
				I29x <= 3039;
				I30x <= 3014;
				I31x <= 3096;
				I32x <= 3153;
				I33x <= 3137;
				I34x <= 2973;
				I35x <= 2777;
				I36x <= 2523;
				I37x <= 2269;
				I38x <= 2056;
				I39x <= 1949;
				I40x <= 1843;
				I41x <= 1720;
				I42x <= 1769;
				I43x <= 1712;
				I44x <= 1777;
				I45x <= 1769;
				I46x <= 1826;
				I47x <= 1843;
				I48x <= 1859;
				I49x <= 1875;
				I50x <= 1933;
				I51x <= 1884;
				I52x <= 1859;
				I53x <= 1810;
				I54x <= 1810;
				I55x <= 1802;
				I56x <= 1744;
				I57x <= 1769;
				I58x <= 1712;
				I59x <= 1720;
				I60x <= 1720;
				I61x <= 1712;
				I62x <= 1785;
				I63x <= 1761;
				I64x <= 1794;
				I65x <= 1802;
				I66x <= 1802;
				I67x <= 1851;
				I68x <= 1859;
				I69x <= 1851;
				I70x <= 1892;
				I71x <= 1884;
				I72x <= 1875;
				I73x <= 1875;
				I74x <= 1859;
				I75x <= 1843;
				I76x <= 1949;
				I77x <= 2113;
				I78x <= 2277;
				I79x <= 2605;
				I80x <= 2850;
				I81x <= 2899;
				I82x <= 2908;
				I83x <= 2383;
				I84x <= 2220;
				I85x <= 2179;
				I86x <= 1933;
				I87x <= 1679;
				I88x <= 1605;
				I89x <= 1712;
				I90x <= 1662;
				I91x <= 1703;
				I92x <= 1736;
				I93x <= 1687;
				I94x <= 1753;
				I95x <= 1802;
				I96x <= 1843;
				I97x <= 1843;
				I98x <= 2179;
				I99x <= 2588;
				I100x <= 3817;
				I101x <= 6717;
				I102x <= 8192;
				I103x <= 3694;
				I104x <= 2211;
				I105x <= 860;
				I106x <= 1048;
				I107x <= 1859;
				I108x <= 2293;
				I109x <= 2359;
				I110x <= 2400;
				I111x <= 2367;
				I112x <= 2490;
				I113x <= 2531;
				I114x <= 2523;
				I115x <= 2629;
				I116x <= 2646;
				I117x <= 2686;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001100:begin
				I0x <= 8192;
				I1x <= 6946;
				I2x <= 2981;
				I3x <= 1392;
				I4x <= 0;
				I5x <= 1114;
				I6x <= 2252;
				I7x <= 2375;
				I8x <= 2523;
				I9x <= 2719;
				I10x <= 2760;
				I11x <= 2859;
				I12x <= 2924;
				I13x <= 2940;
				I14x <= 2883;
				I15x <= 2949;
				I16x <= 3006;
				I17x <= 3039;
				I18x <= 3153;
				I19x <= 3145;
				I20x <= 3153;
				I21x <= 3203;
				I22x <= 3342;
				I23x <= 3391;
				I24x <= 3530;
				I25x <= 3760;
				I26x <= 3956;
				I27x <= 4243;
				I28x <= 4579;
				I29x <= 4849;
				I30x <= 5111;
				I31x <= 5431;
				I32x <= 5545;
				I33x <= 5627;
				I34x <= 5734;
				I35x <= 5603;
				I36x <= 5373;
				I37x <= 4890;
				I38x <= 4399;
				I39x <= 3833;
				I40x <= 3399;
				I41x <= 3096;
				I42x <= 2916;
				I43x <= 2760;
				I44x <= 2719;
				I45x <= 2605;
				I46x <= 2646;
				I47x <= 2596;
				I48x <= 2514;
				I49x <= 2514;
				I50x <= 2506;
				I51x <= 2473;
				I52x <= 2514;
				I53x <= 2580;
				I54x <= 2564;
				I55x <= 2580;
				I56x <= 2580;
				I57x <= 2572;
				I58x <= 2596;
				I59x <= 2605;
				I60x <= 2572;
				I61x <= 2605;
				I62x <= 2605;
				I63x <= 2605;
				I64x <= 2588;
				I65x <= 2539;
				I66x <= 2531;
				I67x <= 2482;
				I68x <= 2473;
				I69x <= 2555;
				I70x <= 2514;
				I71x <= 2441;
				I72x <= 2473;
				I73x <= 2433;
				I74x <= 2457;
				I75x <= 2473;
				I76x <= 2424;
				I77x <= 2408;
				I78x <= 2367;
				I79x <= 2433;
				I80x <= 2424;
				I81x <= 2433;
				I82x <= 2433;
				I83x <= 2457;
				I84x <= 2457;
				I85x <= 2449;
				I86x <= 2400;
				I87x <= 2367;
				I88x <= 2424;
				I89x <= 2408;
				I90x <= 2433;
				I91x <= 2408;
				I92x <= 2424;
				I93x <= 2465;
				I94x <= 2416;
				I95x <= 2441;
				I96x <= 2457;
				I97x <= 2473;
				I98x <= 2473;
				I99x <= 2392;
				I100x <= 2449;
				I101x <= 2490;
				I102x <= 2564;
				I103x <= 2711;
				I104x <= 2727;
				I105x <= 2924;
				I106x <= 2908;
				I107x <= 2818;
				I108x <= 2572;
				I109x <= 2719;
				I110x <= 2555;
				I111x <= 2785;
				I112x <= 2629;
				I113x <= 2531;
				I114x <= 2367;
				I115x <= 2465;
				I116x <= 2498;
				I117x <= 2555;
				I118x <= 2514;
				I119x <= 2596;
				I120x <= 2629;
				I121x <= 2686;
				I122x <= 3039;
				I123x <= 3989;
				I124x <= 4407;
				I125x <= 5931;
				I126x <= 7880;
				I127x <= 5914;
				I128x <= 3121;
				I129x <= 1564;
				I130x <= 516;
				I131x <= 1884;
				I132x <= 2768;
				I133x <= 2801;
				I134x <= 2990;
				I135x <= 3162;
				I136x <= 3252;
				I137x <= 3317;
				I138x <= 3342;
				I139x <= 3383;
				I140x <= 3465;
				I141x <= 3424;
				I142x <= 3489;
				I143x <= 3579;
				I144x <= 3596;
				I145x <= 3661;
				I146x <= 3686;
				I147x <= 3768;
				I148x <= 3850;
				I149x <= 3956;
				I150x <= 4120;
				I151x <= 4284;
				I152x <= 4521;
				I153x <= 4751;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001101:begin
				I0x <= 8192;
				I1x <= 4636;
				I2x <= 1818;
				I3x <= 79;
				I4x <= 262;
				I5x <= 942;
				I6x <= 1384;
				I7x <= 1613;
				I8x <= 1679;
				I9x <= 1753;
				I10x <= 1802;
				I11x <= 1769;
				I12x <= 1720;
				I13x <= 1744;
				I14x <= 1810;
				I15x <= 1810;
				I16x <= 1843;
				I17x <= 1884;
				I18x <= 1908;
				I19x <= 1966;
				I20x <= 2007;
				I21x <= 2080;
				I22x <= 2146;
				I23x <= 2162;
				I24x <= 2318;
				I25x <= 2416;
				I26x <= 2596;
				I27x <= 2744;
				I28x <= 2883;
				I29x <= 3006;
				I30x <= 3162;
				I31x <= 3252;
				I32x <= 3284;
				I33x <= 3153;
				I34x <= 2990;
				I35x <= 2662;
				I36x <= 2482;
				I37x <= 2301;
				I38x <= 2179;
				I39x <= 2031;
				I40x <= 1949;
				I41x <= 1875;
				I42x <= 1867;
				I43x <= 1851;
				I44x <= 1851;
				I45x <= 1794;
				I46x <= 1859;
				I47x <= 1859;
				I48x <= 1802;
				I49x <= 1777;
				I50x <= 1794;
				I51x <= 1810;
				I52x <= 1794;
				I53x <= 1810;
				I54x <= 1728;
				I55x <= 1794;
				I56x <= 1728;
				I57x <= 1818;
				I58x <= 1761;
				I59x <= 1826;
				I60x <= 1810;
				I61x <= 1810;
				I62x <= 1785;
				I63x <= 1744;
				I64x <= 1687;
				I65x <= 1630;
				I66x <= 1662;
				I67x <= 1679;
				I68x <= 1712;
				I69x <= 1744;
				I70x <= 1867;
				I71x <= 2023;
				I72x <= 2220;
				I73x <= 2211;
				I74x <= 2301;
				I75x <= 2334;
				I76x <= 2195;
				I77x <= 2236;
				I78x <= 2031;
				I79x <= 1916;
				I80x <= 1736;
				I81x <= 1630;
				I82x <= 1540;
				I83x <= 1507;
				I84x <= 1482;
				I85x <= 1433;
				I86x <= 1433;
				I87x <= 1286;
				I88x <= 974;
				I89x <= 2359;
				I90x <= 4726;
				I91x <= 7553;
				I92x <= 5070;
				I93x <= 2318;
				I94x <= 62;
				I95x <= 0;
				I96x <= 525;
				I97x <= 1228;
				I98x <= 1400;
				I99x <= 1540;
				I100x <= 1540;
				I101x <= 1597;
				I102x <= 1695;
				I103x <= 1703;
				I104x <= 1794;
				I105x <= 1744;
				I106x <= 1794;
				I107x <= 1884;
				I108x <= 1966;
				I109x <= 2023;
				I110x <= 2031;
				I111x <= 2080;
				I112x <= 2097;
				I113x <= 2105;
				I114x <= 2236;
				I115x <= 2318;
				I116x <= 2473;
				I117x <= 2686;
				I118x <= 2809;
				I119x <= 2924;
				I120x <= 2957;
				I121x <= 3219;
				I122x <= 3276;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001110:begin
				I0x <= 8142;
				I1x <= 6840;
				I2x <= 1163;
				I3x <= 63;
				I4x <= 0;
				I5x <= 485;
				I6x <= 1048;
				I7x <= 1130;
				I8x <= 1146;
				I9x <= 1163;
				I10x <= 1187;
				I11x <= 1228;
				I12x <= 1245;
				I13x <= 1269;
				I14x <= 1327;
				I15x <= 1359;
				I16x <= 1368;
				I17x <= 1376;
				I18x <= 1327;
				I19x <= 1417;
				I20x <= 1482;
				I21x <= 1490;
				I22x <= 1515;
				I23x <= 1605;
				I24x <= 1703;
				I25x <= 1818;
				I26x <= 1925;
				I27x <= 2023;
				I28x <= 2138;
				I29x <= 2293;
				I30x <= 2433;
				I31x <= 2629;
				I32x <= 2719;
				I33x <= 2785;
				I34x <= 2727;
				I35x <= 2588;
				I36x <= 2310;
				I37x <= 2064;
				I38x <= 1933;
				I39x <= 1687;
				I40x <= 1630;
				I41x <= 1556;
				I42x <= 1515;
				I43x <= 1482;
				I44x <= 1458;
				I45x <= 1441;
				I46x <= 1507;
				I47x <= 1507;
				I48x <= 1474;
				I49x <= 1490;
				I50x <= 1490;
				I51x <= 1482;
				I52x <= 1507;
				I53x <= 1458;
				I54x <= 1531;
				I55x <= 1548;
				I56x <= 1515;
				I57x <= 1540;
				I58x <= 1515;
				I59x <= 1531;
				I60x <= 1490;
				I61x <= 1490;
				I62x <= 1449;
				I63x <= 1425;
				I64x <= 1433;
				I65x <= 1392;
				I66x <= 1409;
				I67x <= 1343;
				I68x <= 1343;
				I69x <= 1392;
				I70x <= 1392;
				I71x <= 1359;
				I72x <= 1376;
				I73x <= 1368;
				I74x <= 1384;
				I75x <= 1376;
				I76x <= 1433;
				I77x <= 1597;
				I78x <= 1957;
				I79x <= 1933;
				I80x <= 1835;
				I81x <= 2228;
				I82x <= 2383;
				I83x <= 2310;
				I84x <= 2252;
				I85x <= 2072;
				I86x <= 1859;
				I87x <= 1613;
				I88x <= 1400;
				I89x <= 1146;
				I90x <= 1130;
				I91x <= 1097;
				I92x <= 1081;
				I93x <= 1015;
				I94x <= 991;
				I95x <= 1024;
				I96x <= 1015;
				I97x <= 652;
				I98x <= 950;
				I99x <= 3309;
				I100x <= 5963;
				I101x <= 7405;
				I102x <= 8192;
				I103x <= 3014;
				I104x <= 207;
				I105x <= 39;
				I106x <= 370;
				I107x <= 779;
				I108x <= 1146;
				I109x <= 1130;
				I110x <= 1130;
				I111x <= 1179;
				I112x <= 1196;
				I113x <= 1196;
				I114x <= 1236;
				I115x <= 1261;
				I116x <= 1277;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00001111:begin
				I0x <= 7831;
				I1x <= 4849;
				I2x <= 1081;
				I3x <= 1097;
				I4x <= 1605;
				I5x <= 3317;
				I6x <= 2883;
				I7x <= 2433;
				I8x <= 2654;
				I9x <= 2514;
				I10x <= 2523;
				I11x <= 2662;
				I12x <= 2744;
				I13x <= 2809;
				I14x <= 2768;
				I15x <= 2981;
				I16x <= 3088;
				I17x <= 3194;
				I18x <= 3465;
				I19x <= 3571;
				I20x <= 3923;
				I21x <= 3981;
				I22x <= 4268;
				I23x <= 4513;
				I24x <= 4767;
				I25x <= 5079;
				I26x <= 5275;
				I27x <= 5341;
				I28x <= 5480;
				I29x <= 5464;
				I30x <= 5480;
				I31x <= 5373;
				I32x <= 5218;
				I33x <= 4980;
				I34x <= 4374;
				I35x <= 4055;
				I36x <= 3579;
				I37x <= 3465;
				I38x <= 3514;
				I39x <= 3121;
				I40x <= 3268;
				I41x <= 3137;
				I42x <= 3104;
				I43x <= 3162;
				I44x <= 3080;
				I45x <= 3047;
				I46x <= 2957;
				I47x <= 3014;
				I48x <= 3252;
				I49x <= 3039;
				I50x <= 3112;
				I51x <= 3096;
				I52x <= 2916;
				I53x <= 3260;
				I54x <= 3014;
				I55x <= 3047;
				I56x <= 2760;
				I57x <= 2940;
				I58x <= 3309;
				I59x <= 3358;
				I60x <= 3842;
				I61x <= 3997;
				I62x <= 4358;
				I63x <= 4456;
				I64x <= 4669;
				I65x <= 4669;
				I66x <= 4890;
				I67x <= 4718;
				I68x <= 4251;
				I69x <= 3809;
				I70x <= 3260;
				I71x <= 2908;
				I72x <= 2457;
				I73x <= 2646;
				I74x <= 2514;
				I75x <= 2539;
				I76x <= 2400;
				I77x <= 2179;
				I78x <= 2547;
				I79x <= 3006;
				I80x <= 4489;
				I81x <= 8192;
				I82x <= 7700;
				I83x <= 4308;
				I84x <= 0;
				I85x <= 1310;
				I86x <= 2203;
				I87x <= 3629;
				I88x <= 2973;
				I89x <= 2596;
				I90x <= 2605;
				I91x <= 2605;
				I92x <= 2605;
				I93x <= 2793;
				I94x <= 2637;
				I95x <= 3047;
				I96x <= 2908;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010000:begin
				I0x <= 8110;
				I1x <= 7831;
				I2x <= 3719;
				I3x <= 618;
				I4x <= 0;
				I5x <= 208;
				I6x <= 498;
				I7x <= 444;
				I8x <= 392;
				I9x <= 456;
				I10x <= 520;
				I11x <= 627;
				I12x <= 589;
				I13x <= 708;
				I14x <= 755;
				I15x <= 776;
				I16x <= 851;
				I17x <= 991;
				I18x <= 1097;
				I19x <= 1187;
				I20x <= 1302;
				I21x <= 1572;
				I22x <= 1826;
				I23x <= 2007;
				I24x <= 2220;
				I25x <= 2588;
				I26x <= 2965;
				I27x <= 3203;
				I28x <= 3563;
				I29x <= 3678;
				I30x <= 3891;
				I31x <= 3973;
				I32x <= 3842;
				I33x <= 3383;
				I34x <= 2785;
				I35x <= 2252;
				I36x <= 1810;
				I37x <= 1384;
				I38x <= 1015;
				I39x <= 801;
				I40x <= 529;
				I41x <= 606;
				I42x <= 563;
				I43x <= 550;
				I44x <= 507;
				I45x <= 550;
				I46x <= 541;
				I47x <= 486;
				I48x <= 520;
				I49x <= 494;
				I50x <= 601;
				I51x <= 652;
				I52x <= 639;
				I53x <= 635;
				I54x <= 712;
				I55x <= 724;
				I56x <= 597;
				I57x <= 601;
				I58x <= 665;
				I59x <= 670;
				I60x <= 597;
				I61x <= 584;
				I62x <= 610;
				I63x <= 550;
				I64x <= 503;
				I65x <= 533;
				I66x <= 494;
				I67x <= 486;
				I68x <= 512;
				I69x <= 460;
				I70x <= 512;
				I71x <= 426;
				I72x <= 503;
				I73x <= 520;
				I74x <= 507;
				I75x <= 498;
				I76x <= 439;
				I77x <= 482;
				I78x <= 448;
				I79x <= 434;
				I80x <= 541;
				I81x <= 665;
				I82x <= 876;
				I83x <= 835;
				I84x <= 815;
				I85x <= 1196;
				I86x <= 1310;
				I87x <= 1097;
				I88x <= 884;
				I89x <= 901;
				I90x <= 703;
				I91x <= 486;
				I92x <= 388;
				I93x <= 324;
				I94x <= 303;
				I95x <= 299;
				I96x <= 299;
				I97x <= 230;
				I98x <= 264;
				I99x <= 264;
				I100x <= 149;
				I101x <= 763;
				I102x <= 1425;
				I103x <= 4104;
				I104x <= 8192;
				I105x <= 7831;
				I106x <= 4268;
				I107x <= 909;
				I108x <= 63;
				I109x <= 332;
				I110x <= 554;
				I111x <= 631;
				I112x <= 537;
				I113x <= 656;
				I114x <= 546;
				I115x <= 695;
				I116x <= 665;
				I117x <= 815;
				I118x <= 851;
				I119x <= 933;
				I120x <= 983;
				I121x <= 1130;
				I122x <= 1130;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010001:begin
				I0x <= 7544;
				I1x <= 5578;
				I2x <= 1441;
				I3x <= 884;
				I4x <= 1163;
				I5x <= 1499;
				I6x <= 1499;
				I7x <= 1458;
				I8x <= 1474;
				I9x <= 1327;
				I10x <= 1359;
				I11x <= 1253;
				I12x <= 1220;
				I13x <= 1212;
				I14x <= 1212;
				I15x <= 1327;
				I16x <= 1376;
				I17x <= 1441;
				I18x <= 1458;
				I19x <= 1548;
				I20x <= 1818;
				I21x <= 1794;
				I22x <= 1966;
				I23x <= 2220;
				I24x <= 2531;
				I25x <= 2719;
				I26x <= 3072;
				I27x <= 3440;
				I28x <= 3522;
				I29x <= 3973;
				I30x <= 4186;
				I31x <= 4005;
				I32x <= 3497;
				I33x <= 3235;
				I34x <= 2793;
				I35x <= 2252;
				I36x <= 1941;
				I37x <= 1597;
				I38x <= 1114;
				I39x <= 1163;
				I40x <= 901;
				I41x <= 835;
				I42x <= 724;
				I43x <= 933;
				I44x <= 1187;
				I45x <= 1007;
				I46x <= 958;
				I47x <= 1130;
				I48x <= 1105;
				I49x <= 1146;
				I50x <= 1073;
				I51x <= 1327;
				I52x <= 1212;
				I53x <= 1286;
				I54x <= 1196;
				I55x <= 1064;
				I56x <= 884;
				I57x <= 1007;
				I58x <= 1048;
				I59x <= 1073;
				I60x <= 1048;
				I61x <= 983;
				I62x <= 1163;
				I63x <= 983;
				I64x <= 763;
				I65x <= 851;
				I66x <= 860;
				I67x <= 768;
				I68x <= 753;
				I69x <= 699;
				I70x <= 813;
				I71x <= 589;
				I72x <= 884;
				I73x <= 1220;
				I74x <= 1114;
				I75x <= 1679;
				I76x <= 2105;
				I77x <= 2228;
				I78x <= 2228;
				I79x <= 1720;
				I80x <= 1474;
				I81x <= 788;
				I82x <= 516;
				I83x <= 490;
				I84x <= 321;
				I85x <= 188;
				I86x <= 0;
				I87x <= 44;
				I88x <= 173;
				I89x <= 69;
				I90x <= 625;
				I91x <= 2441;
				I92x <= 4694;
				I93x <= 8192;
				I94x <= 5177;
				I95x <= 1073;
				I96x <= 421;
				I97x <= 892;
				I98x <= 1466;
				I99x <= 1351;
				I100x <= 1327;
				I101x <= 1368;
				I102x <= 1286;
				I103x <= 1638;
				I104x <= 1245;
				I105x <= 1449;
				I106x <= 1302;
				I107x <= 1490;
				I108x <= 1490;
				I109x <= 1466;
				I110x <= 1392;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010010:begin
				I0x <= 7749;
				I1x <= 7651;
				I2x <= 5292;
				I3x <= 2375;
				I4x <= 575;
				I5x <= 0;
				I6x <= 424;
				I7x <= 800;
				I8x <= 776;
				I9x <= 788;
				I10x <= 800;
				I11x <= 814;
				I12x <= 851;
				I13x <= 876;
				I14x <= 950;
				I15x <= 974;
				I16x <= 991;
				I17x <= 1015;
				I18x <= 1056;
				I19x <= 1056;
				I20x <= 1122;
				I21x <= 1220;
				I22x <= 1318;
				I23x <= 1384;
				I24x <= 1433;
				I25x <= 1556;
				I26x <= 1654;
				I27x <= 1810;
				I28x <= 1966;
				I29x <= 2170;
				I30x <= 2359;
				I31x <= 2564;
				I32x <= 2727;
				I33x <= 2834;
				I34x <= 2949;
				I35x <= 2965;
				I36x <= 2940;
				I37x <= 2875;
				I38x <= 2662;
				I39x <= 2375;
				I40x <= 2097;
				I41x <= 1826;
				I42x <= 1597;
				I43x <= 1351;
				I44x <= 1212;
				I45x <= 1097;
				I46x <= 1015;
				I47x <= 933;
				I48x <= 925;
				I49x <= 950;
				I50x <= 942;
				I51x <= 901;
				I52x <= 925;
				I53x <= 933;
				I54x <= 950;
				I55x <= 958;
				I56x <= 925;
				I57x <= 950;
				I58x <= 942;
				I59x <= 958;
				I60x <= 950;
				I61x <= 909;
				I62x <= 950;
				I63x <= 917;
				I64x <= 909;
				I65x <= 950;
				I66x <= 933;
				I67x <= 917;
				I68x <= 892;
				I69x <= 876;
				I70x <= 851;
				I71x <= 819;
				I72x <= 835;
				I73x <= 811;
				I74x <= 797;
				I75x <= 788;
				I76x <= 800;
				I77x <= 791;
				I78x <= 768;
				I79x <= 761;
				I80x <= 802;
				I81x <= 770;
				I82x <= 776;
				I83x <= 756;
				I84x <= 802;
				I85x <= 800;
				I86x <= 759;
				I87x <= 750;
				I88x <= 733;
				I89x <= 756;
				I90x <= 768;
				I91x <= 791;
				I92x <= 779;
				I93x <= 715;
				I94x <= 727;
				I95x <= 759;
				I96x <= 776;
				I97x <= 774;
				I98x <= 802;
				I99x <= 782;
				I100x <= 827;
				I101x <= 793;
				I102x <= 802;
				I103x <= 782;
				I104x <= 793;
				I105x <= 782;
				I106x <= 851;
				I107x <= 999;
				I108x <= 1228;
				I109x <= 1392;
				I110x <= 1597;
				I111x <= 1736;
				I112x <= 1859;
				I113x <= 1843;
				I114x <= 1728;
				I115x <= 1515;
				I116x <= 1441;
				I117x <= 1261;
				I118x <= 901;
				I119x <= 709;
				I120x <= 663;
				I121x <= 628;
				I122x <= 639;
				I123x <= 645;
				I124x <= 599;
				I125x <= 343;
				I126x <= 611;
				I127x <= 2236;
				I128x <= 5865;
				I129x <= 8192;
				I130x <= 7462;
				I131x <= 3964;
				I132x <= 1818;
				I133x <= 194;
				I134x <= 369;
				I135x <= 942;
				I136x <= 966;
				I137x <= 925;
				I138x <= 974;
				I139x <= 1032;
				I140x <= 1040;
				I141x <= 1064;
				I142x <= 1097;
				I143x <= 1105;
				I144x <= 1171;
				I145x <= 1220;
				I146x <= 1286;
				I147x <= 1286;
				I148x <= 1351;
				I149x <= 1433;
				I150x <= 1482;
				I151x <= 1499;
				I152x <= 1622;
				I153x <= 1728;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010011:begin
				I0x <= 7839;
				I1x <= 5660;
				I2x <= 2981;
				I3x <= 1261;
				I4x <= 484;
				I5x <= 1810;
				I6x <= 2465;
				I7x <= 2547;
				I8x <= 2678;
				I9x <= 2875;
				I10x <= 2940;
				I11x <= 2908;
				I12x <= 3022;
				I13x <= 3088;
				I14x <= 3162;
				I15x <= 3121;
				I16x <= 3178;
				I17x <= 3325;
				I18x <= 3358;
				I19x <= 3465;
				I20x <= 3473;
				I21x <= 3596;
				I22x <= 3702;
				I23x <= 3899;
				I24x <= 4153;
				I25x <= 4505;
				I26x <= 4743;
				I27x <= 4915;
				I28x <= 5038;
				I29x <= 5242;
				I30x <= 5349;
				I31x <= 5382;
				I32x <= 5242;
				I33x <= 5005;
				I34x <= 4579;
				I35x <= 4194;
				I36x <= 3776;
				I37x <= 3489;
				I38x <= 3252;
				I39x <= 3039;
				I40x <= 2908;
				I41x <= 2883;
				I42x <= 2891;
				I43x <= 2793;
				I44x <= 2752;
				I45x <= 2736;
				I46x <= 2809;
				I47x <= 2768;
				I48x <= 2744;
				I49x <= 2785;
				I50x <= 2768;
				I51x <= 2834;
				I52x <= 2744;
				I53x <= 2801;
				I54x <= 2883;
				I55x <= 2842;
				I56x <= 2785;
				I57x <= 2785;
				I58x <= 2850;
				I59x <= 2752;
				I60x <= 2686;
				I61x <= 2711;
				I62x <= 2678;
				I63x <= 2621;
				I64x <= 2686;
				I65x <= 2670;
				I66x <= 2629;
				I67x <= 2621;
				I68x <= 2572;
				I69x <= 2637;
				I70x <= 2588;
				I71x <= 2547;
				I72x <= 2482;
				I73x <= 2441;
				I74x <= 2465;
				I75x <= 2408;
				I76x <= 2408;
				I77x <= 2449;
				I78x <= 2433;
				I79x <= 2433;
				I80x <= 2433;
				I81x <= 2490;
				I82x <= 2449;
				I83x <= 2465;
				I84x <= 2400;
				I85x <= 2400;
				I86x <= 2424;
				I87x <= 2506;
				I88x <= 2777;
				I89x <= 3039;
				I90x <= 3088;
				I91x <= 3375;
				I92x <= 3645;
				I93x <= 3497;
				I94x <= 3424;
				I95x <= 3457;
				I96x <= 3129;
				I97x <= 2867;
				I98x <= 2555;
				I99x <= 2318;
				I100x <= 2285;
				I101x <= 2310;
				I102x <= 2269;
				I103x <= 2392;
				I104x <= 2334;
				I105x <= 2252;
				I106x <= 2301;
				I107x <= 2662;
				I108x <= 3563;
				I109x <= 3973;
				I110x <= 5480;
				I111x <= 8192;
				I112x <= 6643;
				I113x <= 3260;
				I114x <= 1032;
				I115x <= 0;
				I116x <= 1376;
				I117x <= 2236;
				I118x <= 2375;
				I119x <= 2572;
				I120x <= 2768;
				I121x <= 2777;
				I122x <= 2752;
				I123x <= 2850;
				I124x <= 2826;
				I125x <= 2965;
				I126x <= 3031;
				I127x <= 3047;
				I128x <= 3104;
				I129x <= 3203;
				I130x <= 3325;
				I131x <= 3440;
				I132x <= 3579;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010100:begin
				I0x <= 8192;
				I1x <= 4341;
				I2x <= 1875;
				I3x <= 868;
				I4x <= 1130;
				I5x <= 2162;
				I6x <= 2310;
				I7x <= 2580;
				I8x <= 2678;
				I9x <= 2883;
				I10x <= 2908;
				I11x <= 2965;
				I12x <= 2965;
				I13x <= 2899;
				I14x <= 2891;
				I15x <= 2990;
				I16x <= 2990;
				I17x <= 3055;
				I18x <= 3006;
				I19x <= 2957;
				I20x <= 3031;
				I21x <= 3088;
				I22x <= 3031;
				I23x <= 3145;
				I24x <= 3358;
				I25x <= 3440;
				I26x <= 3465;
				I27x <= 3440;
				I28x <= 3678;
				I29x <= 3833;
				I30x <= 3907;
				I31x <= 4177;
				I32x <= 4415;
				I33x <= 4644;
				I34x <= 4907;
				I35x <= 4956;
				I36x <= 5120;
				I37x <= 5144;
				I38x <= 5038;
				I39x <= 4841;
				I40x <= 4513;
				I41x <= 4145;
				I42x <= 3883;
				I43x <= 3588;
				I44x <= 3342;
				I45x <= 3055;
				I46x <= 3022;
				I47x <= 2916;
				I48x <= 2818;
				I49x <= 2875;
				I50x <= 2899;
				I51x <= 2940;
				I52x <= 3055;
				I53x <= 2990;
				I54x <= 2998;
				I55x <= 3006;
				I56x <= 3170;
				I57x <= 3162;
				I58x <= 3080;
				I59x <= 3096;
				I60x <= 2998;
				I61x <= 3022;
				I62x <= 2998;
				I63x <= 2965;
				I64x <= 3031;
				I65x <= 2859;
				I66x <= 2859;
				I67x <= 2809;
				I68x <= 2809;
				I69x <= 2752;
				I70x <= 2670;
				I71x <= 2678;
				I72x <= 2678;
				I73x <= 2605;
				I74x <= 2564;
				I75x <= 2555;
				I76x <= 2613;
				I77x <= 2564;
				I78x <= 2473;
				I79x <= 2506;
				I80x <= 2465;
				I81x <= 2457;
				I82x <= 2424;
				I83x <= 2334;
				I84x <= 2293;
				I85x <= 2334;
				I86x <= 2392;
				I87x <= 2408;
				I88x <= 2334;
				I89x <= 2351;
				I90x <= 2301;
				I91x <= 2408;
				I92x <= 2326;
				I93x <= 2310;
				I94x <= 2326;
				I95x <= 2342;
				I96x <= 2490;
				I97x <= 2629;
				I98x <= 2621;
				I99x <= 2727;
				I100x <= 2957;
				I101x <= 2998;
				I102x <= 2670;
				I103x <= 2408;
				I104x <= 2228;
				I105x <= 2072;
				I106x <= 2015;
				I107x <= 1900;
				I108x <= 1892;
				I109x <= 1843;
				I110x <= 1884;
				I111x <= 1941;
				I112x <= 1990;
				I113x <= 1925;
				I114x <= 1892;
				I115x <= 1851;
				I116x <= 1794;
				I117x <= 1720;
				I118x <= 1949;
				I119x <= 2621;
				I120x <= 2924;
				I121x <= 5431;
				I122x <= 7725;
				I123x <= 3637;
				I124x <= 819;
				I125x <= 0;
				I126x <= 530;
				I127x <= 1548;
				I128x <= 1638;
				I129x <= 1818;
				I130x <= 2007;
				I131x <= 2170;
				I132x <= 2236;
				I133x <= 2195;
				I134x <= 2260;
				I135x <= 2342;
				I136x <= 2351;
				I137x <= 2392;
				I138x <= 2334;
				I139x <= 2383;
				I140x <= 2416;
				I141x <= 2457;
				I142x <= 2473;
				I143x <= 2490;
				I144x <= 2580;
				I145x <= 2605;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010101:begin
				I0x <= 7946;
				I1x <= 1957;
				I2x <= 98;
				I3x <= 0;
				I4x <= 1122;
				I5x <= 1310;
				I6x <= 1310;
				I7x <= 1138;
				I8x <= 1138;
				I9x <= 1220;
				I10x <= 1171;
				I11x <= 1212;
				I12x <= 1212;
				I13x <= 1204;
				I14x <= 1351;
				I15x <= 1286;
				I16x <= 1351;
				I17x <= 1409;
				I18x <= 1466;
				I19x <= 1589;
				I20x <= 1671;
				I21x <= 1671;
				I22x <= 1736;
				I23x <= 1802;
				I24x <= 1875;
				I25x <= 2015;
				I26x <= 2195;
				I27x <= 2342;
				I28x <= 2531;
				I29x <= 2703;
				I30x <= 2883;
				I31x <= 3039;
				I32x <= 3178;
				I33x <= 3391;
				I34x <= 3514;
				I35x <= 3629;
				I36x <= 3735;
				I37x <= 3670;
				I38x <= 3563;
				I39x <= 3309;
				I40x <= 3055;
				I41x <= 2768;
				I42x <= 2490;
				I43x <= 2277;
				I44x <= 2187;
				I45x <= 2113;
				I46x <= 2048;
				I47x <= 2007;
				I48x <= 1925;
				I49x <= 1933;
				I50x <= 1925;
				I51x <= 1949;
				I52x <= 1900;
				I53x <= 1892;
				I54x <= 1826;
				I55x <= 1826;
				I56x <= 1835;
				I57x <= 1802;
				I58x <= 1818;
				I59x <= 1810;
				I60x <= 1818;
				I61x <= 1802;
				I62x <= 1810;
				I63x <= 1818;
				I64x <= 1892;
				I65x <= 1794;
				I66x <= 1843;
				I67x <= 1761;
				I68x <= 1794;
				I69x <= 1744;
				I70x <= 1695;
				I71x <= 1777;
				I72x <= 1777;
				I73x <= 1703;
				I74x <= 1753;
				I75x <= 1720;
				I76x <= 1703;
				I77x <= 1695;
				I78x <= 1753;
				I79x <= 1662;
				I80x <= 1695;
				I81x <= 1769;
				I82x <= 1695;
				I83x <= 1900;
				I84x <= 2162;
				I85x <= 2269;
				I86x <= 2220;
				I87x <= 2359;
				I88x <= 2367;
				I89x <= 2228;
				I90x <= 2367;
				I91x <= 2408;
				I92x <= 2293;
				I93x <= 2252;
				I94x <= 2170;
				I95x <= 2097;
				I96x <= 1744;
				I97x <= 1556;
				I98x <= 1589;
				I99x <= 1630;
				I100x <= 1482;
				I101x <= 1466;
				I102x <= 1581;
				I103x <= 1523;
				I104x <= 1515;
				I105x <= 1482;
				I106x <= 1982;
				I107x <= 2940;
				I108x <= 5144;
				I109x <= 6758;
				I110x <= 8192;
				I111x <= 2383;
				I112x <= 494;
				I113x <= 253;
				I114x <= 1286;
				I115x <= 1572;
				I116x <= 1597;
				I117x <= 1458;
				I118x <= 1474;
				I119x <= 1499;
				I120x <= 1507;
				I121x <= 1531;
				I122x <= 1507;
				I123x <= 1466;
				I124x <= 1531;
				I125x <= 1581;
				I126x <= 1613;
				I127x <= 1630;
				I128x <= 1744;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010110:begin
				I0x <= 7806;
				I1x <= 4571;
				I2x <= 1990;
				I3x <= 767;
				I4x <= 983;
				I5x <= 835;
				I6x <= 733;
				I7x <= 706;
				I8x <= 475;
				I9x <= 706;
				I10x <= 654;
				I11x <= 514;
				I12x <= 662;
				I13x <= 475;
				I14x <= 697;
				I15x <= 645;
				I16x <= 610;
				I17x <= 763;
				I18x <= 649;
				I19x <= 909;
				I20x <= 901;
				I21x <= 860;
				I22x <= 942;
				I23x <= 724;
				I24x <= 1040;
				I25x <= 999;
				I26x <= 1040;
				I27x <= 1261;
				I28x <= 1163;
				I29x <= 1482;
				I30x <= 1466;
				I31x <= 1490;
				I32x <= 1826;
				I33x <= 1720;
				I34x <= 2056;
				I35x <= 2154;
				I36x <= 2162;
				I37x <= 2400;
				I38x <= 2056;
				I39x <= 2121;
				I40x <= 1859;
				I41x <= 1679;
				I42x <= 1695;
				I43x <= 1253;
				I44x <= 1286;
				I45x <= 983;
				I46x <= 876;
				I47x <= 983;
				I48x <= 763;
				I49x <= 974;
				I50x <= 966;
				I51x <= 933;
				I52x <= 933;
				I53x <= 645;
				I54x <= 901;
				I55x <= 950;
				I56x <= 860;
				I57x <= 925;
				I58x <= 711;
				I59x <= 815;
				I60x <= 715;
				I61x <= 589;
				I62x <= 693;
				I63x <= 488;
				I64x <= 784;
				I65x <= 733;
				I66x <= 680;
				I67x <= 827;
				I68x <= 584;
				I69x <= 793;
				I70x <= 759;
				I71x <= 619;
				I72x <= 662;
				I73x <= 440;
				I74x <= 771;
				I75x <= 602;
				I76x <= 532;
				I77x <= 641;
				I78x <= 466;
				I79x <= 606;
				I80x <= 789;
				I81x <= 658;
				I82x <= 750;
				I83x <= 558;
				I84x <= 675;
				I85x <= 545;
				I86x <= 606;
				I87x <= 759;
				I88x <= 497;
				I89x <= 684;
				I90x <= 733;
				I91x <= 680;
				I92x <= 827;
				I93x <= 553;
				I94x <= 702;
				I95x <= 693;
				I96x <= 671;
				I97x <= 649;
				I98x <= 435;
				I99x <= 806;
				I100x <= 767;
				I101x <= 759;
				I102x <= 884;
				I103x <= 706;
				I104x <= 868;
				I105x <= 892;
				I106x <= 759;
				I107x <= 860;
				I108x <= 632;
				I109x <= 950;
				I110x <= 1097;
				I111x <= 1466;
				I112x <= 1515;
				I113x <= 1302;
				I114x <= 1572;
				I115x <= 1736;
				I116x <= 1351;
				I117x <= 1318;
				I118x <= 860;
				I119x <= 1097;
				I120x <= 1122;
				I121x <= 811;
				I122x <= 835;
				I123x <= 510;
				I124x <= 784;
				I125x <= 724;
				I126x <= 667;
				I127x <= 645;
				I128x <= 0;
				I129x <= 1024;
				I130x <= 4014;
				I131x <= 6807;
				I132x <= 8192;
				I133x <= 4620;
				I134x <= 1933;
				I135x <= 733;
				I136x <= 793;
				I137x <= 784;
				I138x <= 532;
				I139x <= 641;
				I140x <= 597;
				I141x <= 545;
				I142x <= 584;
				I143x <= 484;
				I144x <= 549;
				I145x <= 602;
				I146x <= 558;
				I147x <= 793;
				I148x <= 584;
				I149x <= 715;
				I150x <= 675;
				I151x <= 649;
				I152x <= 901;
				I153x <= 593;
				I154x <= 917;
				I155x <= 835;
				I156x <= 827;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00010111:begin
				I0x <= 8192;
				I1x <= 5644;
				I2x <= 3407;
				I3x <= 384;
				I4x <= 137;
				I5x <= 1146;
				I6x <= 1851;
				I7x <= 2154;
				I8x <= 2113;
				I9x <= 2252;
				I10x <= 2260;
				I11x <= 2236;
				I12x <= 2424;
				I13x <= 2351;
				I14x <= 2457;
				I15x <= 2433;
				I16x <= 2400;
				I17x <= 2564;
				I18x <= 2457;
				I19x <= 2621;
				I20x <= 2547;
				I21x <= 2506;
				I22x <= 2662;
				I23x <= 2572;
				I24x <= 2711;
				I25x <= 2711;
				I26x <= 2727;
				I27x <= 2981;
				I28x <= 3055;
				I29x <= 3162;
				I30x <= 2940;
				I31x <= 2678;
				I32x <= 2629;
				I33x <= 2367;
				I34x <= 2285;
				I35x <= 2203;
				I36x <= 2244;
				I37x <= 2228;
				I38x <= 2039;
				I39x <= 2121;
				I40x <= 2121;
				I41x <= 2015;
				I42x <= 2203;
				I43x <= 2121;
				I44x <= 2203;
				I45x <= 2236;
				I46x <= 2228;
				I47x <= 2555;
				I48x <= 2752;
				I49x <= 2940;
				I50x <= 3031;
				I51x <= 3153;
				I52x <= 3252;
				I53x <= 3317;
				I54x <= 3375;
				I55x <= 3186;
				I56x <= 2859;
				I57x <= 2564;
				I58x <= 2138;
				I59x <= 2088;
				I60x <= 1957;
				I61x <= 1777;
				I62x <= 1884;
				I63x <= 1761;
				I64x <= 1802;
				I65x <= 1736;
				I66x <= 1654;
				I67x <= 1744;
				I68x <= 1548;
				I69x <= 1974;
				I70x <= 2662;
				I71x <= 5701;
				I72x <= 7716;
				I73x <= 4489;
				I74x <= 2678;
				I75x <= 0;
				I76x <= 144;
				I77x <= 1236;
				I78x <= 1802;
				I79x <= 1957;
				I80x <= 1966;
				I81x <= 1941;
				I82x <= 2105;
				I83x <= 2056;
				I84x <= 2179;
				I85x <= 0;
				I86x <= 0;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011000:begin
				I0x <= 8192;
				I1x <= 6029;
				I2x <= 2285;
				I3x <= 702;
				I4x <= 1220;
				I5x <= 1196;
				I6x <= 1024;
				I7x <= 1015;
				I8x <= 1007;
				I9x <= 942;
				I10x <= 983;
				I11x <= 983;
				I12x <= 1048;
				I13x <= 1114;
				I14x <= 1138;
				I15x <= 1105;
				I16x <= 1187;
				I17x <= 1089;
				I18x <= 1212;
				I19x <= 1196;
				I20x <= 1277;
				I21x <= 1277;
				I22x <= 1277;
				I23x <= 1433;
				I24x <= 1523;
				I25x <= 1482;
				I26x <= 1597;
				I27x <= 1703;
				I28x <= 1916;
				I29x <= 2064;
				I30x <= 2203;
				I31x <= 2433;
				I32x <= 2744;
				I33x <= 3129;
				I34x <= 3276;
				I35x <= 3481;
				I36x <= 3514;
				I37x <= 3432;
				I38x <= 3088;
				I39x <= 2703;
				I40x <= 2318;
				I41x <= 1875;
				I42x <= 1728;
				I43x <= 1400;
				I44x <= 1228;
				I45x <= 1179;
				I46x <= 1122;
				I47x <= 892;
				I48x <= 1015;
				I49x <= 942;
				I50x <= 809;
				I51x <= 933;
				I52x <= 868;
				I53x <= 787;
				I54x <= 884;
				I55x <= 925;
				I56x <= 892;
				I57x <= 868;
				I58x <= 860;
				I59x <= 909;
				I60x <= 991;
				I61x <= 974;
				I62x <= 1007;
				I63x <= 966;
				I64x <= 974;
				I65x <= 958;
				I66x <= 925;
				I67x <= 819;
				I68x <= 764;
				I69x <= 819;
				I70x <= 773;
				I71x <= 715;
				I72x <= 729;
				I73x <= 729;
				I74x <= 706;
				I75x <= 764;
				I76x <= 711;
				I77x <= 800;
				I78x <= 778;
				I79x <= 738;
				I80x <= 634;
				I81x <= 760;
				I82x <= 773;
				I83x <= 729;
				I84x <= 742;
				I85x <= 711;
				I86x <= 764;
				I87x <= 715;
				I88x <= 679;
				I89x <= 720;
				I90x <= 751;
				I91x <= 738;
				I92x <= 652;
				I93x <= 697;
				I94x <= 693;
				I95x <= 819;
				I96x <= 1048;
				I97x <= 1212;
				I98x <= 1359;
				I99x <= 1261;
				I100x <= 1212;
				I101x <= 1466;
				I102x <= 1392;
				I103x <= 1171;
				I104x <= 1097;
				I105x <= 917;
				I106x <= 796;
				I107x <= 742;
				I108x <= 634;
				I109x <= 536;
				I110x <= 625;
				I111x <= 576;
				I112x <= 581;
				I113x <= 518;
				I114x <= 598;
				I115x <= 523;
				I116x <= 67;
				I117x <= 0;
				I118x <= 1531;
				I119x <= 6127;
				I120x <= 8110;
				I121x <= 6201;
				I122x <= 2252;
				I123x <= 549;
				I124x <= 1056;
				I125x <= 1089;
				I126x <= 884;
				I127x <= 892;
				I128x <= 851;
				I129x <= 909;
				I130x <= 925;
				I131x <= 909;
				I132x <= 860;
				I133x <= 958;
				I134x <= 958;
				I135x <= 983;
				I136x <= 942;
				I137x <= 999;
				I138x <= 1089;
				I139x <= 1146;
				I140x <= 1253;
				I141x <= 1212;
				I142x <= 1228;
				I143x <= 1302;
				I144x <= 1351;
				I145x <= 1400;
				I146x <= 1482;
				I147x <= 1523;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011001:begin
				I0x <= 8192;
				I1x <= 6578;
				I2x <= 2629;
				I3x <= 534;
				I4x <= 1703;
				I5x <= 3031;
				I6x <= 3342;
				I7x <= 2899;
				I8x <= 2654;
				I9x <= 2834;
				I10x <= 2932;
				I11x <= 2719;
				I12x <= 2801;
				I13x <= 2957;
				I14x <= 3014;
				I15x <= 3104;
				I16x <= 3162;
				I17x <= 3301;
				I18x <= 3334;
				I19x <= 3547;
				I20x <= 3612;
				I21x <= 3710;
				I22x <= 4005;
				I23x <= 4104;
				I24x <= 4333;
				I25x <= 4644;
				I26x <= 4595;
				I27x <= 4947;
				I28x <= 4816;
				I29x <= 4849;
				I30x <= 5021;
				I31x <= 4825;
				I32x <= 4792;
				I33x <= 4530;
				I34x <= 4349;
				I35x <= 3997;
				I36x <= 3563;
				I37x <= 3383;
				I38x <= 3178;
				I39x <= 3137;
				I40x <= 3203;
				I41x <= 2981;
				I42x <= 2998;
				I43x <= 2850;
				I44x <= 3096;
				I45x <= 3153;
				I46x <= 2990;
				I47x <= 3088;
				I48x <= 2998;
				I49x <= 3121;
				I50x <= 3072;
				I51x <= 2768;
				I52x <= 2973;
				I53x <= 2899;
				I54x <= 2932;
				I55x <= 3244;
				I56x <= 3293;
				I57x <= 3702;
				I58x <= 3858;
				I59x <= 4005;
				I60x <= 4259;
				I61x <= 4145;
				I62x <= 4292;
				I63x <= 4366;
				I64x <= 4153;
				I65x <= 3751;
				I66x <= 3203;
				I67x <= 2867;
				I68x <= 2621;
				I69x <= 2473;
				I70x <= 2383;
				I71x <= 2334;
				I72x <= 2244;
				I73x <= 2236;
				I74x <= 2285;
				I75x <= 2678;
				I76x <= 2785;
				I77x <= 4603;
				I78x <= 7471;
				I79x <= 5709;
				I80x <= 1908;
				I81x <= 0;
				I82x <= 1040;
				I83x <= 2621;
				I84x <= 2875;
				I85x <= 2367;
				I86x <= 2203;
				I87x <= 2236;
				I88x <= 2334;
				I89x <= 2392;
				I90x <= 2506;
				I91x <= 2621;
				I92x <= 2637;
				I93x <= 2654;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011010:begin
				I0x <= 7716;
				I1x <= 6602;
				I2x <= 3506;
				I3x <= 1523;
				I4x <= 186;
				I5x <= 600;
				I6x <= 1146;
				I7x <= 1146;
				I8x <= 1171;
				I9x <= 1155;
				I10x <= 1196;
				I11x <= 1179;
				I12x <= 1204;
				I13x <= 1204;
				I14x <= 1220;
				I15x <= 1220;
				I16x <= 1236;
				I17x <= 1269;
				I18x <= 1351;
				I19x <= 1376;
				I20x <= 1409;
				I21x <= 1433;
				I22x <= 1548;
				I23x <= 1654;
				I24x <= 1753;
				I25x <= 1851;
				I26x <= 1957;
				I27x <= 2072;
				I28x <= 2170;
				I29x <= 2228;
				I30x <= 2252;
				I31x <= 2326;
				I32x <= 2277;
				I33x <= 2301;
				I34x <= 2072;
				I35x <= 1867;
				I36x <= 1646;
				I37x <= 1441;
				I38x <= 1269;
				I39x <= 1130;
				I40x <= 1032;
				I41x <= 983;
				I42x <= 925;
				I43x <= 925;
				I44x <= 884;
				I45x <= 909;
				I46x <= 974;
				I47x <= 901;
				I48x <= 974;
				I49x <= 958;
				I50x <= 991;
				I51x <= 1024;
				I52x <= 991;
				I53x <= 999;
				I54x <= 1007;
				I55x <= 1024;
				I56x <= 991;
				I57x <= 966;
				I58x <= 999;
				I59x <= 925;
				I60x <= 892;
				I61x <= 876;
				I62x <= 851;
				I63x <= 851;
				I64x <= 799;
				I65x <= 799;
				I66x <= 797;
				I67x <= 753;
				I68x <= 747;
				I69x <= 741;
				I70x <= 711;
				I71x <= 735;
				I72x <= 670;
				I73x <= 686;
				I74x <= 677;
				I75x <= 704;
				I76x <= 720;
				I77x <= 714;
				I78x <= 711;
				I79x <= 674;
				I80x <= 686;
				I81x <= 695;
				I82x <= 670;
				I83x <= 707;
				I84x <= 677;
				I85x <= 738;
				I86x <= 753;
				I87x <= 692;
				I88x <= 738;
				I89x <= 892;
				I90x <= 1081;
				I91x <= 1032;
				I92x <= 942;
				I93x <= 868;
				I94x <= 772;
				I95x <= 763;
				I96x <= 760;
				I97x <= 707;
				I98x <= 677;
				I99x <= 517;
				I100x <= 410;
				I101x <= 438;
				I102x <= 420;
				I103x <= 480;
				I104x <= 456;
				I105x <= 487;
				I106x <= 557;
				I107x <= 551;
				I108x <= 607;
				I109x <= 554;
				I110x <= 621;
				I111x <= 1744;
				I112x <= 5226;
				I113x <= 8192;
				I114x <= 4472;
				I115x <= 2555;
				I116x <= 524;
				I117x <= 0;
				I118x <= 536;
				I119x <= 950;
				I120x <= 884;
				I121x <= 819;
				I122x <= 892;
				I123x <= 876;
				I124x <= 942;
				I125x <= 925;
				I126x <= 983;
				I127x <= 950;
				I128x <= 991;
				I129x <= 999;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011011:begin
				I0x <= 7995;
				I1x <= 7905;
				I2x <= 3244;
				I3x <= 966;
				I4x <= 623;
				I5x <= 1671;
				I6x <= 2318;
				I7x <= 2613;
				I8x <= 2703;
				I9x <= 2703;
				I10x <= 2760;
				I11x <= 2801;
				I12x <= 2826;
				I13x <= 2793;
				I14x <= 2826;
				I15x <= 2826;
				I16x <= 2867;
				I17x <= 2899;
				I18x <= 2842;
				I19x <= 2883;
				I20x <= 2957;
				I21x <= 3047;
				I22x <= 3104;
				I23x <= 3211;
				I24x <= 3407;
				I25x <= 3620;
				I26x <= 3809;
				I27x <= 4030;
				I28x <= 4284;
				I29x <= 4513;
				I30x <= 4767;
				I31x <= 4923;
				I32x <= 5013;
				I33x <= 5070;
				I34x <= 4997;
				I35x <= 4784;
				I36x <= 4431;
				I37x <= 4022;
				I38x <= 3588;
				I39x <= 3211;
				I40x <= 2908;
				I41x <= 2777;
				I42x <= 2596;
				I43x <= 2523;
				I44x <= 2392;
				I45x <= 2293;
				I46x <= 2277;
				I47x <= 2211;
				I48x <= 2170;
				I49x <= 2179;
				I50x <= 2195;
				I51x <= 2228;
				I52x <= 2301;
				I53x <= 2342;
				I54x <= 2351;
				I55x <= 2342;
				I56x <= 2351;
				I57x <= 2375;
				I58x <= 2375;
				I59x <= 2293;
				I60x <= 2285;
				I61x <= 2244;
				I62x <= 2211;
				I63x <= 2211;
				I64x <= 2244;
				I65x <= 2260;
				I66x <= 2244;
				I67x <= 2195;
				I68x <= 2138;
				I69x <= 2064;
				I70x <= 1982;
				I71x <= 1941;
				I72x <= 1941;
				I73x <= 1949;
				I74x <= 1908;
				I75x <= 1867;
				I76x <= 1843;
				I77x <= 1859;
				I78x <= 1933;
				I79x <= 1908;
				I80x <= 1949;
				I81x <= 1998;
				I82x <= 1892;
				I83x <= 1859;
				I84x <= 1843;
				I85x <= 1859;
				I86x <= 1867;
				I87x <= 1900;
				I88x <= 1908;
				I89x <= 1908;
				I90x <= 1966;
				I91x <= 1982;
				I92x <= 1957;
				I93x <= 1949;
				I94x <= 1916;
				I95x <= 1933;
				I96x <= 1933;
				I97x <= 2031;
				I98x <= 2105;
				I99x <= 2113;
				I100x <= 2170;
				I101x <= 2146;
				I102x <= 2146;
				I103x <= 2424;
				I104x <= 2646;
				I105x <= 2457;
				I106x <= 2359;
				I107x <= 2031;
				I108x <= 1982;
				I109x <= 1908;
				I110x <= 1925;
				I111x <= 1900;
				I112x <= 1908;
				I113x <= 1900;
				I114x <= 1916;
				I115x <= 1916;
				I116x <= 1925;
				I117x <= 1941;
				I118x <= 1884;
				I119x <= 1818;
				I120x <= 1785;
				I121x <= 2580;
				I122x <= 4153;
				I123x <= 5971;
				I124x <= 8192;
				I125x <= 5070;
				I126x <= 1400;
				I127x <= 0;
				I128x <= 752;
				I129x <= 1622;
				I130x <= 2039;
				I131x <= 2121;
				I132x <= 2113;
				I133x <= 2097;
				I134x <= 2154;
				I135x <= 2146;
				I136x <= 2211;
				I137x <= 2236;
				I138x <= 2269;
				I139x <= 2301;
				I140x <= 2334;
				I141x <= 2367;
				I142x <= 2441;
				I143x <= 2572;
				I144x <= 2629;
				I145x <= 2711;
				I146x <= 2809;
				I147x <= 2957;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011100:begin
				I0x <= 8101;
				I1x <= 6504;
				I2x <= 3923;
				I3x <= 2048;
				I4x <= 1359;
				I5x <= 1605;
				I6x <= 1679;
				I7x <= 1622;
				I8x <= 1613;
				I9x <= 1622;
				I10x <= 1646;
				I11x <= 1679;
				I12x <= 1671;
				I13x <= 1679;
				I14x <= 1687;
				I15x <= 1744;
				I16x <= 1777;
				I17x <= 1826;
				I18x <= 1875;
				I19x <= 1925;
				I20x <= 2015;
				I21x <= 2088;
				I22x <= 2195;
				I23x <= 2301;
				I24x <= 2416;
				I25x <= 2555;
				I26x <= 2686;
				I27x <= 2768;
				I28x <= 2859;
				I29x <= 2908;
				I30x <= 2957;
				I31x <= 2981;
				I32x <= 2850;
				I33x <= 2670;
				I34x <= 2449;
				I35x <= 2220;
				I36x <= 2039;
				I37x <= 1884;
				I38x <= 1761;
				I39x <= 1703;
				I40x <= 1646;
				I41x <= 1646;
				I42x <= 1662;
				I43x <= 1662;
				I44x <= 1638;
				I45x <= 1630;
				I46x <= 1654;
				I47x <= 1622;
				I48x <= 1662;
				I49x <= 1671;
				I50x <= 1662;
				I51x <= 1671;
				I52x <= 1646;
				I53x <= 1662;
				I54x <= 1654;
				I55x <= 1671;
				I56x <= 1671;
				I57x <= 1662;
				I58x <= 1630;
				I59x <= 1720;
				I60x <= 1802;
				I61x <= 1892;
				I62x <= 1941;
				I63x <= 1990;
				I64x <= 2129;
				I65x <= 2203;
				I66x <= 2244;
				I67x <= 2203;
				I68x <= 2039;
				I69x <= 1761;
				I70x <= 1564;
				I71x <= 1515;
				I72x <= 1449;
				I73x <= 1458;
				I74x <= 1417;
				I75x <= 1441;
				I76x <= 1425;
				I77x <= 1466;
				I78x <= 1433;
				I79x <= 1449;
				I80x <= 1441;
				I81x <= 1449;
				I82x <= 1155;
				I83x <= 0;
				I84x <= 835;
				I85x <= 2990;
				I86x <= 6021;
				I87x <= 8192;
				I88x <= 5079;
				I89x <= 3317;
				I90x <= 1622;
				I91x <= 1531;
				I92x <= 1794;
				I93x <= 1843;
				I94x <= 1794;
				I95x <= 1777;
				I96x <= 1785;
				I97x <= 1802;
				I98x <= 1826;
				I99x <= 1859;
				I100x <= 1859;
				I101x <= 1900;
				I102x <= 1957;
				I103x <= 2007;
				I104x <= 2056;
				I105x <= 2113;
				I106x <= 2211;
				I107x <= 2334;
				I108x <= 2408;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011101:begin
				I0x <= 7888;
				I1x <= 8192;
				I2x <= 2375;
				I3x <= 638;
				I4x <= 337;
				I5x <= 476;
				I6x <= 1220;
				I7x <= 1490;
				I8x <= 1458;
				I9x <= 1490;
				I10x <= 1482;
				I11x <= 1515;
				I12x <= 1540;
				I13x <= 1589;
				I14x <= 1687;
				I15x <= 1703;
				I16x <= 1777;
				I17x <= 1802;
				I18x <= 1794;
				I19x <= 1761;
				I20x <= 1859;
				I21x <= 1908;
				I22x <= 2007;
				I23x <= 2088;
				I24x <= 2203;
				I25x <= 2310;
				I26x <= 2424;
				I27x <= 2506;
				I28x <= 2613;
				I29x <= 2760;
				I30x <= 2990;
				I31x <= 3276;
				I32x <= 3489;
				I33x <= 3702;
				I34x <= 3915;
				I35x <= 4128;
				I36x <= 4284;
				I37x <= 4349;
				I38x <= 4317;
				I39x <= 4087;
				I40x <= 3694;
				I41x <= 3284;
				I42x <= 2859;
				I43x <= 2473;
				I44x <= 2129;
				I45x <= 1916;
				I46x <= 1687;
				I47x <= 1564;
				I48x <= 1466;
				I49x <= 1392;
				I50x <= 1351;
				I51x <= 1327;
				I52x <= 1351;
				I53x <= 1343;
				I54x <= 1351;
				I55x <= 1425;
				I56x <= 1400;
				I57x <= 1449;
				I58x <= 1417;
				I59x <= 1433;
				I60x <= 1507;
				I61x <= 1540;
				I62x <= 1605;
				I63x <= 1613;
				I64x <= 1581;
				I65x <= 1540;
				I66x <= 1441;
				I67x <= 1376;
				I68x <= 1392;
				I69x <= 1376;
				I70x <= 1327;
				I71x <= 1351;
				I72x <= 1310;
				I73x <= 1318;
				I74x <= 1318;
				I75x <= 1286;
				I76x <= 1245;
				I77x <= 1261;
				I78x <= 1286;
				I79x <= 1286;
				I80x <= 1220;
				I81x <= 1236;
				I82x <= 1228;
				I83x <= 1179;
				I84x <= 1196;
				I85x <= 1220;
				I86x <= 1204;
				I87x <= 1138;
				I88x <= 1089;
				I89x <= 1179;
				I90x <= 1138;
				I91x <= 1155;
				I92x <= 1097;
				I93x <= 1114;
				I94x <= 1081;
				I95x <= 1089;
				I96x <= 1105;
				I97x <= 1122;
				I98x <= 1089;
				I99x <= 1081;
				I100x <= 1081;
				I101x <= 1048;
				I102x <= 1097;
				I103x <= 1122;
				I104x <= 1179;
				I105x <= 1515;
				I106x <= 1671;
				I107x <= 1794;
				I108x <= 1843;
				I109x <= 1966;
				I110x <= 1933;
				I111x <= 1769;
				I112x <= 1556;
				I113x <= 1376;
				I114x <= 1286;
				I115x <= 1081;
				I116x <= 933;
				I117x <= 925;
				I118x <= 884;
				I119x <= 843;
				I120x <= 806;
				I121x <= 788;
				I122x <= 762;
				I123x <= 795;
				I124x <= 747;
				I125x <= 362;
				I126x <= 868;
				I127x <= 4194;
				I128x <= 7741;
				I129x <= 7380;
				I130x <= 1671;
				I131x <= 245;
				I132x <= 0;
				I133x <= 282;
				I134x <= 983;
				I135x <= 1146;
				I136x <= 1155;
				I137x <= 1179;
				I138x <= 1171;
				I139x <= 1179;
				I140x <= 1212;
				I141x <= 1269;
				I142x <= 1261;
				I143x <= 1277;
				I144x <= 1294;
				I145x <= 1368;
				I146x <= 1400;
				I147x <= 1384;
				I148x <= 1409;
				I149x <= 1482;
				I150x <= 1589;
				I151x <= 1662;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011110:begin
				I0x <= 8192;
				I1x <= 4096;
				I2x <= 715;
				I3x <= 513;
				I4x <= 1204;
				I5x <= 1564;
				I6x <= 1810;
				I7x <= 1875;
				I8x <= 1867;
				I9x <= 1941;
				I10x <= 2097;
				I11x <= 2007;
				I12x <= 1982;
				I13x <= 1949;
				I14x <= 2228;
				I15x <= 2048;
				I16x <= 2252;
				I17x <= 2097;
				I18x <= 2154;
				I19x <= 2269;
				I20x <= 2408;
				I21x <= 2473;
				I22x <= 2473;
				I23x <= 2736;
				I24x <= 2809;
				I25x <= 2940;
				I26x <= 3112;
				I27x <= 3457;
				I28x <= 3530;
				I29x <= 3760;
				I30x <= 3874;
				I31x <= 3891;
				I32x <= 3932;
				I33x <= 3842;
				I34x <= 3563;
				I35x <= 3309;
				I36x <= 3055;
				I37x <= 2686;
				I38x <= 2678;
				I39x <= 2367;
				I40x <= 2269;
				I41x <= 2154;
				I42x <= 2293;
				I43x <= 2195;
				I44x <= 2097;
				I45x <= 2220;
				I46x <= 2113;
				I47x <= 2228;
				I48x <= 2252;
				I49x <= 2162;
				I50x <= 2351;
				I51x <= 2375;
				I52x <= 2277;
				I53x <= 2334;
				I54x <= 2359;
				I55x <= 2228;
				I56x <= 2228;
				I57x <= 2326;
				I58x <= 2129;
				I59x <= 2146;
				I60x <= 2105;
				I61x <= 1998;
				I62x <= 2097;
				I63x <= 2015;
				I64x <= 2154;
				I65x <= 1974;
				I66x <= 2072;
				I67x <= 2187;
				I68x <= 2031;
				I69x <= 2015;
				I70x <= 2121;
				I71x <= 2277;
				I72x <= 2482;
				I73x <= 2760;
				I74x <= 2908;
				I75x <= 2981;
				I76x <= 2695;
				I77x <= 2981;
				I78x <= 2646;
				I79x <= 2310;
				I80x <= 2203;
				I81x <= 2154;
				I82x <= 1908;
				I83x <= 2064;
				I84x <= 1867;
				I85x <= 1777;
				I86x <= 1867;
				I87x <= 1826;
				I88x <= 1769;
				I89x <= 1679;
				I90x <= 1785;
				I91x <= 1662;
				I92x <= 1687;
				I93x <= 1220;
				I94x <= 1581;
				I95x <= 3588;
				I96x <= 4931;
				I97x <= 7036;
				I98x <= 5398;
				I99x <= 1458;
				I100x <= 0;
				I101x <= 561;
				I102x <= 1155;
				I103x <= 1531;
				I104x <= 1777;
				I105x <= 1818;
				I106x <= 1769;
				I107x <= 1916;
				I108x <= 1818;
				I109x <= 1843;
				I110x <= 1949;
				I111x <= 1998;
				I112x <= 1966;
				I113x <= 1867;
				I114x <= 1998;
				I115x <= 2080;
				I116x <= 2064;
				I117x <= 2236;
				I118x <= 2514;
				I119x <= 2506;
				I120x <= 2506;
				I121x <= 2572;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00011111:begin
				I0x <= 7340;
				I1x <= 7536;
				I2x <= 3866;
				I3x <= 2015;
				I4x <= 404;
				I5x <= 699;
				I6x <= 2072;
				I7x <= 2441;
				I8x <= 2580;
				I9x <= 2736;
				I10x <= 2801;
				I11x <= 2908;
				I12x <= 2973;
				I13x <= 3047;
				I14x <= 3039;
				I15x <= 3006;
				I16x <= 3080;
				I17x <= 3178;
				I18x <= 3186;
				I19x <= 3244;
				I20x <= 3440;
				I21x <= 3497;
				I22x <= 3670;
				I23x <= 3825;
				I24x <= 4145;
				I25x <= 4374;
				I26x <= 4743;
				I27x <= 5079;
				I28x <= 5242;
				I29x <= 5414;
				I30x <= 5529;
				I31x <= 5521;
				I32x <= 5242;
				I33x <= 4808;
				I34x <= 4349;
				I35x <= 3784;
				I36x <= 3309;
				I37x <= 3022;
				I38x <= 2727;
				I39x <= 2596;
				I40x <= 2605;
				I41x <= 2539;
				I42x <= 2441;
				I43x <= 2416;
				I44x <= 2375;
				I45x <= 2433;
				I46x <= 2367;
				I47x <= 2359;
				I48x <= 2326;
				I49x <= 2342;
				I50x <= 2310;
				I51x <= 2285;
				I52x <= 2351;
				I53x <= 2310;
				I54x <= 2457;
				I55x <= 2441;
				I56x <= 2433;
				I57x <= 2400;
				I58x <= 2326;
				I59x <= 2400;
				I60x <= 2351;
				I61x <= 2392;
				I62x <= 2293;
				I63x <= 2392;
				I64x <= 2334;
				I65x <= 2260;
				I66x <= 2187;
				I67x <= 2236;
				I68x <= 2236;
				I69x <= 2187;
				I70x <= 2203;
				I71x <= 2162;
				I72x <= 2154;
				I73x <= 2138;
				I74x <= 2121;
				I75x <= 2138;
				I76x <= 2187;
				I77x <= 2121;
				I78x <= 2048;
				I79x <= 2105;
				I80x <= 2105;
				I81x <= 2080;
				I82x <= 2064;
				I83x <= 2236;
				I84x <= 2326;
				I85x <= 2457;
				I86x <= 2490;
				I87x <= 2416;
				I88x <= 2383;
				I89x <= 2310;
				I90x <= 2236;
				I91x <= 2400;
				I92x <= 2236;
				I93x <= 2195;
				I94x <= 2064;
				I95x <= 1941;
				I96x <= 2015;
				I97x <= 2080;
				I98x <= 2113;
				I99x <= 2088;
				I100x <= 2146;
				I101x <= 2228;
				I102x <= 2465;
				I103x <= 3407;
				I104x <= 3596;
				I105x <= 5038;
				I106x <= 8192;
				I107x <= 6889;
				I108x <= 3145;
				I109x <= 1122;
				I110x <= 0;
				I111x <= 1261;
				I112x <= 2187;
				I113x <= 2310;
				I114x <= 2596;
				I115x <= 2686;
				I116x <= 2842;
				I117x <= 2867;
				I118x <= 2826;
				I119x <= 2965;
				I120x <= 2916;
				I121x <= 2940;
				I122x <= 3031;
				I123x <= 3080;
				I124x <= 3162;
				I125x <= 3268;
				I126x <= 3301;
				I127x <= 3407;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100000:begin
				I0x <= 8192;
				I1x <= 5308;
				I2x <= 1368;
				I3x <= 813;
				I4x <= 1187;
				I5x <= 1507;
				I6x <= 1376;
				I7x <= 1294;
				I8x <= 1318;
				I9x <= 1318;
				I10x <= 1359;
				I11x <= 1359;
				I12x <= 1327;
				I13x <= 1392;
				I14x <= 1384;
				I15x <= 1351;
				I16x <= 1318;
				I17x <= 1318;
				I18x <= 1384;
				I19x <= 1417;
				I20x <= 1449;
				I21x <= 1507;
				I22x <= 1507;
				I23x <= 1654;
				I24x <= 1671;
				I25x <= 1851;
				I26x <= 1941;
				I27x <= 2023;
				I28x <= 2326;
				I29x <= 2523;
				I30x <= 2793;
				I31x <= 3080;
				I32x <= 3293;
				I33x <= 3629;
				I34x <= 3858;
				I35x <= 4046;
				I36x <= 3956;
				I37x <= 3588;
				I38x <= 3121;
				I39x <= 2564;
				I40x <= 2039;
				I41x <= 1679;
				I42x <= 1392;
				I43x <= 1236;
				I44x <= 1105;
				I45x <= 1056;
				I46x <= 1032;
				I47x <= 983;
				I48x <= 1032;
				I49x <= 1015;
				I50x <= 1056;
				I51x <= 991;
				I52x <= 942;
				I53x <= 1015;
				I54x <= 1032;
				I55x <= 1073;
				I56x <= 1073;
				I57x <= 1105;
				I58x <= 1155;
				I59x <= 1064;
				I60x <= 1081;
				I61x <= 1114;
				I62x <= 1097;
				I63x <= 1122;
				I64x <= 1114;
				I65x <= 1138;
				I66x <= 1089;
				I67x <= 1024;
				I68x <= 1024;
				I69x <= 1007;
				I70x <= 1007;
				I71x <= 991;
				I72x <= 901;
				I73x <= 1048;
				I74x <= 1032;
				I75x <= 958;
				I76x <= 909;
				I77x <= 835;
				I78x <= 901;
				I79x <= 851;
				I80x <= 787;
				I81x <= 819;
				I82x <= 743;
				I83x <= 800;
				I84x <= 819;
				I85x <= 790;
				I86x <= 783;
				I87x <= 868;
				I88x <= 1105;
				I89x <= 1138;
				I90x <= 1163;
				I91x <= 1277;
				I92x <= 1286;
				I93x <= 1327;
				I94x <= 1286;
				I95x <= 1105;
				I96x <= 1040;
				I97x <= 925;
				I98x <= 806;
				I99x <= 727;
				I100x <= 704;
				I101x <= 707;
				I102x <= 632;
				I103x <= 625;
				I104x <= 562;
				I105x <= 559;
				I106x <= 582;
				I107x <= 579;
				I108x <= 684;
				I109x <= 684;
				I110x <= 642;
				I111x <= 516;
				I112x <= 0;
				I113x <= 362;
				I114x <= 1581;
				I115x <= 5095;
				I116x <= 7716;
				I117x <= 5824;
				I118x <= 1630;
				I119x <= 299;
				I120x <= 549;
				I121x <= 1089;
				I122x <= 901;
				I123x <= 860;
				I124x <= 851;
				I125x <= 843;
				I126x <= 851;
				I127x <= 892;
				I128x <= 925;
				I129x <= 876;
				I130x <= 909;
				I131x <= 925;
				I132x <= 925;
				I133x <= 909;
				I134x <= 950;
				I135x <= 950;
				I136x <= 1048;
				I137x <= 1064;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100001:begin
				I0x <= 7847;
				I1x <= 3039;
				I2x <= 446;
				I3x <= 0;
				I4x <= 437;
				I5x <= 1581;
				I6x <= 1712;
				I7x <= 2072;
				I8x <= 2154;
				I9x <= 2392;
				I10x <= 2514;
				I11x <= 2572;
				I12x <= 2564;
				I13x <= 2375;
				I14x <= 2514;
				I15x <= 2613;
				I16x <= 2506;
				I17x <= 2473;
				I18x <= 2523;
				I19x <= 2646;
				I20x <= 2670;
				I21x <= 2744;
				I22x <= 2768;
				I23x <= 2916;
				I24x <= 2981;
				I25x <= 3112;
				I26x <= 3268;
				I27x <= 3448;
				I28x <= 3661;
				I29x <= 3842;
				I30x <= 3956;
				I31x <= 4169;
				I32x <= 4505;
				I33x <= 4595;
				I34x <= 4743;
				I35x <= 4988;
				I36x <= 5005;
				I37x <= 4947;
				I38x <= 4882;
				I39x <= 4734;
				I40x <= 4374;
				I41x <= 3923;
				I42x <= 3768;
				I43x <= 3342;
				I44x <= 3178;
				I45x <= 3211;
				I46x <= 2965;
				I47x <= 2867;
				I48x <= 2859;
				I49x <= 2924;
				I50x <= 2981;
				I51x <= 2891;
				I52x <= 2957;
				I53x <= 3022;
				I54x <= 3047;
				I55x <= 2949;
				I56x <= 3104;
				I57x <= 3121;
				I58x <= 3006;
				I59x <= 3112;
				I60x <= 3055;
				I61x <= 2990;
				I62x <= 3080;
				I63x <= 3039;
				I64x <= 3063;
				I65x <= 3047;
				I66x <= 2940;
				I67x <= 2990;
				I68x <= 3055;
				I69x <= 2981;
				I70x <= 2924;
				I71x <= 2809;
				I72x <= 2867;
				I73x <= 2842;
				I74x <= 2826;
				I75x <= 2768;
				I76x <= 2719;
				I77x <= 2859;
				I78x <= 2686;
				I79x <= 2752;
				I80x <= 2768;
				I81x <= 2777;
				I82x <= 2793;
				I83x <= 2744;
				I84x <= 2793;
				I85x <= 2768;
				I86x <= 2719;
				I87x <= 2719;
				I88x <= 2613;
				I89x <= 2580;
				I90x <= 2473;
				I91x <= 2539;
				I92x <= 2605;
				I93x <= 2826;
				I94x <= 3112;
				I95x <= 3022;
				I96x <= 3235;
				I97x <= 3506;
				I98x <= 3309;
				I99x <= 3235;
				I100x <= 2908;
				I101x <= 2482;
				I102x <= 2457;
				I103x <= 2318;
				I104x <= 2244;
				I105x <= 2318;
				I106x <= 2334;
				I107x <= 2269;
				I108x <= 2277;
				I109x <= 2211;
				I110x <= 2203;
				I111x <= 2228;
				I112x <= 2260;
				I113x <= 2064;
				I114x <= 2023;
				I115x <= 2973;
				I116x <= 3137;
				I117x <= 4104;
				I118x <= 8192;
				I119x <= 7192;
				I120x <= 2547;
				I121x <= 288;
				I122x <= 21;
				I123x <= 1114;
				I124x <= 1843;
				I125x <= 2228;
				I126x <= 2351;
				I127x <= 2490;
				I128x <= 2547;
				I129x <= 2596;
				I130x <= 2605;
				I131x <= 2621;
				I132x <= 2637;
				I133x <= 2703;
				I134x <= 2826;
				I135x <= 2727;
				I136x <= 2818;
				I137x <= 3039;
				I138x <= 3080;
				I139x <= 3194;
				I140x <= 3284;
				I141x <= 3235;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100010:begin
				I0x <= 8085;
				I1x <= 7184;
				I2x <= 2334;
				I3x <= 98;
				I4x <= 261;
				I5x <= 807;
				I6x <= 801;
				I7x <= 739;
				I8x <= 709;
				I9x <= 736;
				I10x <= 719;
				I11x <= 787;
				I12x <= 835;
				I13x <= 892;
				I14x <= 909;
				I15x <= 917;
				I16x <= 933;
				I17x <= 991;
				I18x <= 1024;
				I19x <= 1089;
				I20x <= 1105;
				I21x <= 1187;
				I22x <= 1327;
				I23x <= 1449;
				I24x <= 1515;
				I25x <= 1556;
				I26x <= 1736;
				I27x <= 1818;
				I28x <= 1949;
				I29x <= 2252;
				I30x <= 2457;
				I31x <= 2777;
				I32x <= 3072;
				I33x <= 3366;
				I34x <= 3645;
				I35x <= 3809;
				I36x <= 3915;
				I37x <= 3801;
				I38x <= 3325;
				I39x <= 2793;
				I40x <= 2269;
				I41x <= 1826;
				I42x <= 1425;
				I43x <= 1155;
				I44x <= 1024;
				I45x <= 892;
				I46x <= 868;
				I47x <= 868;
				I48x <= 807;
				I49x <= 868;
				I50x <= 814;
				I51x <= 851;
				I52x <= 835;
				I53x <= 851;
				I54x <= 860;
				I55x <= 797;
				I56x <= 835;
				I57x <= 884;
				I58x <= 860;
				I59x <= 843;
				I60x <= 876;
				I61x <= 925;
				I62x <= 950;
				I63x <= 909;
				I64x <= 917;
				I65x <= 827;
				I66x <= 851;
				I67x <= 817;
				I68x <= 787;
				I69x <= 793;
				I70x <= 753;
				I71x <= 807;
				I72x <= 760;
				I73x <= 685;
				I74x <= 725;
				I75x <= 597;
				I76x <= 624;
				I77x <= 668;
				I78x <= 698;
				I79x <= 760;
				I80x <= 682;
				I81x <= 725;
				I82x <= 725;
				I83x <= 709;
				I84x <= 851;
				I85x <= 1073;
				I86x <= 1155;
				I87x <= 1220;
				I88x <= 1351;
				I89x <= 1417;
				I90x <= 1392;
				I91x <= 1318;
				I92x <= 1155;
				I93x <= 1081;
				I94x <= 999;
				I95x <= 807;
				I96x <= 692;
				I97x <= 631;
				I98x <= 590;
				I99x <= 600;
				I100x <= 560;
				I101x <= 549;
				I102x <= 552;
				I103x <= 584;
				I104x <= 614;
				I105x <= 579;
				I106x <= 603;
				I107x <= 549;
				I108x <= 508;
				I109x <= 326;
				I110x <= 0;
				I111x <= 1220;
				I112x <= 3571;
				I113x <= 8192;
				I114x <= 7643;
				I115x <= 2875;
				I116x <= 451;
				I117x <= 444;
				I118x <= 868;
				I119x <= 999;
				I120x <= 884;
				I121x <= 950;
				I122x <= 950;
				I123x <= 917;
				I124x <= 958;
				I125x <= 851;
				I126x <= 966;
				I127x <= 958;
				I128x <= 991;
				I129x <= 1064;
				I130x <= 1015;
				I131x <= 1089;
				I132x <= 1073;
				I133x <= 1179;
				I134x <= 1204;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100011:begin
				I0x <= 8192;
				I1x <= 5341;
				I2x <= 3244;
				I3x <= 1687;
				I4x <= 1630;
				I5x <= 1794;
				I6x <= 1802;
				I7x <= 1761;
				I8x <= 1769;
				I9x <= 1777;
				I10x <= 1802;
				I11x <= 1802;
				I12x <= 1826;
				I13x <= 1843;
				I14x <= 1859;
				I15x <= 1892;
				I16x <= 1941;
				I17x <= 1966;
				I18x <= 1998;
				I19x <= 2080;
				I20x <= 2138;
				I21x <= 2220;
				I22x <= 2318;
				I23x <= 2392;
				I24x <= 2498;
				I25x <= 2637;
				I26x <= 2752;
				I27x <= 2867;
				I28x <= 2940;
				I29x <= 3014;
				I30x <= 3063;
				I31x <= 3112;
				I32x <= 3047;
				I33x <= 2899;
				I34x <= 2662;
				I35x <= 2433;
				I36x <= 2195;
				I37x <= 2039;
				I38x <= 1892;
				I39x <= 1794;
				I40x <= 1761;
				I41x <= 1712;
				I42x <= 1679;
				I43x <= 1695;
				I44x <= 1695;
				I45x <= 1695;
				I46x <= 1695;
				I47x <= 1720;
				I48x <= 1720;
				I49x <= 1720;
				I50x <= 1712;
				I51x <= 1712;
				I52x <= 1712;
				I53x <= 1720;
				I54x <= 1736;
				I55x <= 1728;
				I56x <= 1728;
				I57x <= 1744;
				I58x <= 1744;
				I59x <= 1753;
				I60x <= 1744;
				I61x <= 1695;
				I62x <= 1712;
				I63x <= 1712;
				I64x <= 1703;
				I65x <= 1671;
				I66x <= 1671;
				I67x <= 1662;
				I68x <= 1654;
				I69x <= 1654;
				I70x <= 1662;
				I71x <= 1654;
				I72x <= 1638;
				I73x <= 1630;
				I74x <= 1646;
				I75x <= 1744;
				I76x <= 1875;
				I77x <= 1900;
				I78x <= 1949;
				I79x <= 1974;
				I80x <= 2056;
				I81x <= 2097;
				I82x <= 2211;
				I83x <= 2072;
				I84x <= 1925;
				I85x <= 1695;
				I86x <= 1622;
				I87x <= 1572;
				I88x <= 1531;
				I89x <= 1523;
				I90x <= 1507;
				I91x <= 1490;
				I92x <= 1490;
				I93x <= 1507;
				I94x <= 1482;
				I95x <= 1490;
				I96x <= 1490;
				I97x <= 1474;
				I98x <= 892;
				I99x <= 0;
				I100x <= 1417;
				I101x <= 3588;
				I102x <= 6569;
				I103x <= 7593;
				I104x <= 4440;
				I105x <= 2744;
				I106x <= 1507;
				I107x <= 1654;
				I108x <= 1785;
				I109x <= 1744;
				I110x <= 1728;
				I111x <= 1728;
				I112x <= 1736;
				I113x <= 1753;
				I114x <= 1794;
				I115x <= 1818;
				I116x <= 1826;
				I117x <= 1851;
				I118x <= 1900;
				I119x <= 1933;
				I120x <= 1982;
				I121x <= 2023;
				I122x <= 2080;
				I123x <= 2146;
				I124x <= 2236;
				I125x <= 2334;
				I126x <= 2449;
				I127x <= 2580;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100100:begin
				I0x <= 8192;
				I1x <= 5529;
				I2x <= 3096;
				I3x <= 1171;
				I4x <= 0;
				I5x <= 453;
				I6x <= 1015;
				I7x <= 1097;
				I8x <= 1114;
				I9x <= 1138;
				I10x <= 1105;
				I11x <= 1146;
				I12x <= 1187;
				I13x <= 1212;
				I14x <= 1212;
				I15x <= 1253;
				I16x <= 1294;
				I17x <= 1327;
				I18x <= 1409;
				I19x <= 1425;
				I20x <= 1449;
				I21x <= 1548;
				I22x <= 1605;
				I23x <= 1736;
				I24x <= 1826;
				I25x <= 1916;
				I26x <= 2015;
				I27x <= 2105;
				I28x <= 2170;
				I29x <= 2211;
				I30x <= 2252;
				I31x <= 2236;
				I32x <= 2260;
				I33x <= 2154;
				I34x <= 2007;
				I35x <= 1810;
				I36x <= 1671;
				I37x <= 1499;
				I38x <= 1368;
				I39x <= 1277;
				I40x <= 1212;
				I41x <= 1187;
				I42x <= 1212;
				I43x <= 1179;
				I44x <= 1171;
				I45x <= 1179;
				I46x <= 1179;
				I47x <= 1163;
				I48x <= 1196;
				I49x <= 1212;
				I50x <= 1196;
				I51x <= 1187;
				I52x <= 1187;
				I53x <= 1179;
				I54x <= 1187;
				I55x <= 1163;
				I56x <= 1171;
				I57x <= 1146;
				I58x <= 1114;
				I59x <= 1138;
				I60x <= 1097;
				I61x <= 1089;
				I62x <= 1081;
				I63x <= 1081;
				I64x <= 1073;
				I65x <= 1040;
				I66x <= 1040;
				I67x <= 1024;
				I68x <= 1048;
				I69x <= 1048;
				I70x <= 1048;
				I71x <= 1032;
				I72x <= 1032;
				I73x <= 1040;
				I74x <= 1032;
				I75x <= 1032;
				I76x <= 1056;
				I77x <= 1163;
				I78x <= 1220;
				I79x <= 1310;
				I80x <= 1417;
				I81x <= 1597;
				I82x <= 1482;
				I83x <= 1433;
				I84x <= 1335;
				I85x <= 1253;
				I86x <= 1155;
				I87x <= 1310;
				I88x <= 1187;
				I89x <= 1056;
				I90x <= 909;
				I91x <= 851;
				I92x <= 860;
				I93x <= 909;
				I94x <= 892;
				I95x <= 909;
				I96x <= 950;
				I97x <= 999;
				I98x <= 1007;
				I99x <= 1032;
				I100x <= 1073;
				I101x <= 766;
				I102x <= 1507;
				I103x <= 3244;
				I104x <= 7151;
				I105x <= 7970;
				I106x <= 4104;
				I107x <= 2113;
				I108x <= 479;
				I109x <= 618;
				I110x <= 1155;
				I111x <= 1376;
				I112x <= 1335;
				I113x <= 1335;
				I114x <= 1368;
				I115x <= 1409;
				I116x <= 1417;
				I117x <= 1433;
				I118x <= 1474;
				I119x <= 1507;
				I120x <= 1548;
				I121x <= 1572;
				I122x <= 1638;
				I123x <= 1671;
				I124x <= 1761;
				I125x <= 1802;
				I126x <= 1875;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100101:begin
				I0x <= 7438;
				I1x <= 6463;
				I2x <= 2711;
				I3x <= 593;
				I4x <= 0;
				I5x <= 677;
				I6x <= 901;
				I7x <= 819;
				I8x <= 674;
				I9x <= 724;
				I10x <= 750;
				I11x <= 785;
				I12x <= 801;
				I13x <= 804;
				I14x <= 835;
				I15x <= 827;
				I16x <= 851;
				I17x <= 901;
				I18x <= 884;
				I19x <= 942;
				I20x <= 1007;
				I21x <= 1056;
				I22x <= 1097;
				I23x <= 1130;
				I24x <= 1196;
				I25x <= 1269;
				I26x <= 1351;
				I27x <= 1433;
				I28x <= 1531;
				I29x <= 1679;
				I30x <= 1851;
				I31x <= 2015;
				I32x <= 2228;
				I33x <= 2465;
				I34x <= 2695;
				I35x <= 2916;
				I36x <= 3129;
				I37x <= 3309;
				I38x <= 3383;
				I39x <= 3334;
				I40x <= 3137;
				I41x <= 2826;
				I42x <= 2465;
				I43x <= 2064;
				I44x <= 1712;
				I45x <= 1449;
				I46x <= 1187;
				I47x <= 1040;
				I48x <= 933;
				I49x <= 807;
				I50x <= 804;
				I51x <= 785;
				I52x <= 785;
				I53x <= 740;
				I54x <= 770;
				I55x <= 750;
				I56x <= 763;
				I57x <= 792;
				I58x <= 788;
				I59x <= 795;
				I60x <= 795;
				I61x <= 827;
				I62x <= 807;
				I63x <= 835;
				I64x <= 801;
				I65x <= 843;
				I66x <= 788;
				I67x <= 782;
				I68x <= 779;
				I69x <= 788;
				I70x <= 801;
				I71x <= 782;
				I72x <= 779;
				I73x <= 785;
				I74x <= 766;
				I75x <= 775;
				I76x <= 747;
				I77x <= 738;
				I78x <= 661;
				I79x <= 674;
				I80x <= 667;
				I81x <= 715;
				I82x <= 645;
				I83x <= 661;
				I84x <= 674;
				I85x <= 683;
				I86x <= 667;
				I87x <= 674;
				I88x <= 664;
				I89x <= 642;
				I90x <= 647;
				I91x <= 661;
				I92x <= 664;
				I93x <= 667;
				I94x <= 677;
				I95x <= 679;
				I96x <= 664;
				I97x <= 677;
				I98x <= 661;
				I99x <= 686;
				I100x <= 679;
				I101x <= 715;
				I102x <= 782;
				I103x <= 884;
				I104x <= 1056;
				I105x <= 1220;
				I106x <= 1253;
				I107x <= 1286;
				I108x <= 1409;
				I109x <= 1466;
				I110x <= 1351;
				I111x <= 1196;
				I112x <= 1073;
				I113x <= 958;
				I114x <= 814;
				I115x <= 689;
				I116x <= 642;
				I117x <= 619;
				I118x <= 603;
				I119x <= 622;
				I120x <= 619;
				I121x <= 610;
				I122x <= 622;
				I123x <= 616;
				I124x <= 651;
				I125x <= 670;
				I126x <= 679;
				I127x <= 686;
				I128x <= 686;
				I129x <= 341;
				I130x <= 217;
				I131x <= 1220;
				I132x <= 3112;
				I133x <= 5726;
				I134x <= 8192;
				I135x <= 5251;
				I136x <= 2285;
				I137x <= 571;
				I138x <= 575;
				I139x <= 1097;
				I140x <= 1261;
				I141x <= 1130;
				I142x <= 1122;
				I143x <= 1114;
				I144x <= 1105;
				I145x <= 1097;
				I146x <= 1105;
				I147x <= 1114;
				I148x <= 1130;
				I149x <= 1179;
				I150x <= 1196;
				I151x <= 1204;
				I152x <= 1245;
				I153x <= 1269;
				I154x <= 1286;
				I155x <= 1327;
				I156x <= 1409;
				I157x <= 1466;
				I158x <= 1515;
				I159x <= 1564;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100110:begin
				I0x <= 8192;
				I1x <= 7643;
				I2x <= 3964;
				I3x <= 1204;
				I4x <= 240;
				I5x <= 1982;
				I6x <= 2629;
				I7x <= 2662;
				I8x <= 2899;
				I9x <= 3006;
				I10x <= 3088;
				I11x <= 3039;
				I12x <= 3112;
				I13x <= 3186;
				I14x <= 3276;
				I15x <= 3391;
				I16x <= 3424;
				I17x <= 3448;
				I18x <= 3538;
				I19x <= 3604;
				I20x <= 3727;
				I21x <= 3915;
				I22x <= 4079;
				I23x <= 4218;
				I24x <= 4521;
				I25x <= 4800;
				I26x <= 5079;
				I27x <= 5431;
				I28x <= 5693;
				I29x <= 6004;
				I30x <= 6283;
				I31x <= 6389;
				I32x <= 6258;
				I33x <= 5971;
				I34x <= 5488;
				I35x <= 4833;
				I36x <= 4235;
				I37x <= 3686;
				I38x <= 3284;
				I39x <= 3055;
				I40x <= 2899;
				I41x <= 2777;
				I42x <= 2752;
				I43x <= 2752;
				I44x <= 2703;
				I45x <= 2686;
				I46x <= 2637;
				I47x <= 2605;
				I48x <= 2539;
				I49x <= 2621;
				I50x <= 2744;
				I51x <= 2678;
				I52x <= 2736;
				I53x <= 2605;
				I54x <= 2727;
				I55x <= 2752;
				I56x <= 2727;
				I57x <= 2760;
				I58x <= 2711;
				I59x <= 2785;
				I60x <= 2727;
				I61x <= 2662;
				I62x <= 2760;
				I63x <= 2703;
				I64x <= 2613;
				I65x <= 2678;
				I66x <= 2686;
				I67x <= 2596;
				I68x <= 2555;
				I69x <= 2580;
				I70x <= 2531;
				I71x <= 2449;
				I72x <= 2490;
				I73x <= 2498;
				I74x <= 2473;
				I75x <= 2473;
				I76x <= 2441;
				I77x <= 2351;
				I78x <= 2457;
				I79x <= 2400;
				I80x <= 2424;
				I81x <= 2400;
				I82x <= 2359;
				I83x <= 2351;
				I84x <= 2318;
				I85x <= 2375;
				I86x <= 2375;
				I87x <= 2359;
				I88x <= 2383;
				I89x <= 2318;
				I90x <= 2285;
				I91x <= 2359;
				I92x <= 2285;
				I93x <= 2301;
				I94x <= 2383;
				I95x <= 2211;
				I96x <= 2203;
				I97x <= 2244;
				I98x <= 2195;
				I99x <= 2301;
				I100x <= 2768;
				I101x <= 2957;
				I102x <= 3112;
				I103x <= 3252;
				I104x <= 3284;
				I105x <= 2998;
				I106x <= 3235;
				I107x <= 2949;
				I108x <= 2490;
				I109x <= 2244;
				I110x <= 1966;
				I111x <= 1925;
				I112x <= 1949;
				I113x <= 2007;
				I114x <= 1933;
				I115x <= 2048;
				I116x <= 2048;
				I117x <= 1933;
				I118x <= 2195;
				I119x <= 3178;
				I120x <= 3301;
				I121x <= 4538;
				I122x <= 7200;
				I123x <= 6496;
				I124x <= 3358;
				I125x <= 1097;
				I126x <= 0;
				I127x <= 1417;
				I128x <= 2260;
				I129x <= 2277;
				I130x <= 2383;
				I131x <= 2539;
				I132x <= 2662;
				I133x <= 2752;
				I134x <= 2793;
				I135x <= 2949;
				I136x <= 2916;
				I137x <= 2965;
				I138x <= 3096;
				I139x <= 3137;
				I140x <= 3211;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00100111:begin
				I0x <= 7520;
				I1x <= 5693;
				I2x <= 2801;
				I3x <= 1212;
				I4x <= 0;
				I5x <= 357;
				I6x <= 983;
				I7x <= 1097;
				I8x <= 1122;
				I9x <= 1196;
				I10x <= 1204;
				I11x <= 1269;
				I12x <= 1351;
				I13x <= 1433;
				I14x <= 1449;
				I15x <= 1572;
				I16x <= 1572;
				I17x <= 1646;
				I18x <= 1703;
				I19x <= 1785;
				I20x <= 1753;
				I21x <= 1794;
				I22x <= 1875;
				I23x <= 1957;
				I24x <= 2048;
				I25x <= 2170;
				I26x <= 2293;
				I27x <= 2482;
				I28x <= 2637;
				I29x <= 2760;
				I30x <= 2932;
				I31x <= 2957;
				I32x <= 3031;
				I33x <= 3129;
				I34x <= 3162;
				I35x <= 3088;
				I36x <= 2908;
				I37x <= 2678;
				I38x <= 2433;
				I39x <= 2179;
				I40x <= 1941;
				I41x <= 1859;
				I42x <= 1744;
				I43x <= 1638;
				I44x <= 1531;
				I45x <= 1507;
				I46x <= 1499;
				I47x <= 1490;
				I48x <= 1499;
				I49x <= 1482;
				I50x <= 1540;
				I51x <= 1654;
				I52x <= 1589;
				I53x <= 1564;
				I54x <= 1531;
				I55x <= 1499;
				I56x <= 1449;
				I57x <= 1359;
				I58x <= 1425;
				I59x <= 1441;
				I60x <= 1466;
				I61x <= 1507;
				I62x <= 1466;
				I63x <= 1433;
				I64x <= 1409;
				I65x <= 1433;
				I66x <= 1449;
				I67x <= 1490;
				I68x <= 1490;
				I69x <= 1507;
				I70x <= 1466;
				I71x <= 1449;
				I72x <= 1433;
				I73x <= 1409;
				I74x <= 1359;
				I75x <= 1368;
				I76x <= 1359;
				I77x <= 1400;
				I78x <= 1392;
				I79x <= 1556;
				I80x <= 1572;
				I81x <= 1687;
				I82x <= 1572;
				I83x <= 1564;
				I84x <= 1548;
				I85x <= 1507;
				I86x <= 1466;
				I87x <= 1474;
				I88x <= 1474;
				I89x <= 1466;
				I90x <= 1441;
				I91x <= 1474;
				I92x <= 1515;
				I93x <= 1556;
				I94x <= 1564;
				I95x <= 1712;
				I96x <= 1908;
				I97x <= 2039;
				I98x <= 2080;
				I99x <= 2342;
				I100x <= 2359;
				I101x <= 2596;
				I102x <= 2646;
				I103x <= 2473;
				I104x <= 2269;
				I105x <= 2187;
				I106x <= 2056;
				I107x <= 1671;
				I108x <= 1433;
				I109x <= 1351;
				I110x <= 1417;
				I111x <= 1400;
				I112x <= 1368;
				I113x <= 1343;
				I114x <= 1040;
				I115x <= 1318;
				I116x <= 2088;
				I117x <= 5136;
				I118x <= 8192;
				I119x <= 7200;
				I120x <= 4202;
				I121x <= 2416;
				I122x <= 892;
				I123x <= 194;
				I124x <= 835;
				I125x <= 1392;
				I126x <= 1433;
				I127x <= 1482;
				I128x <= 1540;
				I129x <= 1605;
				I130x <= 1695;
				I131x <= 1744;
				I132x <= 1875;
				I133x <= 1859;
				I134x <= 1835;
				I135x <= 1843;
				I136x <= 1925;
				I137x <= 1957;
				I138x <= 1982;
				I139x <= 2097;
				I140x <= 2113;
				I141x <= 2187;
				I142x <= 2293;
				I143x <= 2408;
				I144x <= 2498;
				I145x <= 2654;
				I146x <= 2785;
				I147x <= 2834;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101000:begin
				I0x <= 8192;
				I1x <= 4726;
				I2x <= 2998;
				I3x <= 1376;
				I4x <= 1335;
				I5x <= 1548;
				I6x <= 1597;
				I7x <= 1548;
				I8x <= 1531;
				I9x <= 1548;
				I10x <= 1572;
				I11x <= 1589;
				I12x <= 1622;
				I13x <= 1605;
				I14x <= 1662;
				I15x <= 1712;
				I16x <= 1744;
				I17x <= 1794;
				I18x <= 1867;
				I19x <= 1941;
				I20x <= 2031;
				I21x <= 2097;
				I22x <= 2211;
				I23x <= 2334;
				I24x <= 2490;
				I25x <= 2613;
				I26x <= 2744;
				I27x <= 2867;
				I28x <= 2973;
				I29x <= 3031;
				I30x <= 3088;
				I31x <= 3080;
				I32x <= 2949;
				I33x <= 2768;
				I34x <= 2531;
				I35x <= 2260;
				I36x <= 2048;
				I37x <= 1867;
				I38x <= 1761;
				I39x <= 1695;
				I40x <= 1605;
				I41x <= 1613;
				I42x <= 1581;
				I43x <= 1589;
				I44x <= 1572;
				I45x <= 1564;
				I46x <= 1556;
				I47x <= 1572;
				I48x <= 1572;
				I49x <= 1581;
				I50x <= 1572;
				I51x <= 1589;
				I52x <= 1613;
				I53x <= 1605;
				I54x <= 1613;
				I55x <= 1605;
				I56x <= 1622;
				I57x <= 1589;
				I58x <= 1581;
				I59x <= 1589;
				I60x <= 1613;
				I61x <= 1581;
				I62x <= 1556;
				I63x <= 1548;
				I64x <= 1548;
				I65x <= 1523;
				I66x <= 1531;
				I67x <= 1515;
				I68x <= 1507;
				I69x <= 1490;
				I70x <= 1515;
				I71x <= 1482;
				I72x <= 1482;
				I73x <= 1515;
				I74x <= 1630;
				I75x <= 1720;
				I76x <= 1777;
				I77x <= 1753;
				I78x <= 1843;
				I79x <= 1982;
				I80x <= 1982;
				I81x <= 2015;
				I82x <= 1892;
				I83x <= 1662;
				I84x <= 1449;
				I85x <= 1376;
				I86x <= 1310;
				I87x <= 1277;
				I88x <= 1245;
				I89x <= 1236;
				I90x <= 1253;
				I91x <= 1245;
				I92x <= 1236;
				I93x <= 1228;
				I94x <= 1220;
				I95x <= 1228;
				I96x <= 1105;
				I97x <= 49;
				I98x <= 0;
				I99x <= 2080;
				I100x <= 5079;
				I101x <= 8192;
				I102x <= 6078;
				I103x <= 3612;
				I104x <= 1753;
				I105x <= 1253;
				I106x <= 1474;
				I107x <= 1507;
				I108x <= 1458;
				I109x <= 1449;
				I110x <= 1466;
				I111x <= 1482;
				I112x <= 1507;
				I113x <= 1523;
				I114x <= 1540;
				I115x <= 1556;
				I116x <= 1572;
				I117x <= 1613;
				I118x <= 1662;
				I119x <= 1720;
				I120x <= 1769;
				I121x <= 1859;
				I122x <= 1933;
				I123x <= 2031;
				I124x <= 2162;
				I125x <= 2285;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101001:begin
				I0x <= 8192;
				I1x <= 4177;
				I2x <= 416;
				I3x <= 480;
				I4x <= 535;
				I5x <= 465;
				I6x <= 299;
				I7x <= 286;
				I8x <= 286;
				I9x <= 316;
				I10x <= 239;
				I11x <= 217;
				I12x <= 197;
				I13x <= 222;
				I14x <= 250;
				I15x <= 282;
				I16x <= 296;
				I17x <= 270;
				I18x <= 316;
				I19x <= 354;
				I20x <= 385;
				I21x <= 403;
				I22x <= 480;
				I23x <= 561;
				I24x <= 682;
				I25x <= 827;
				I26x <= 991;
				I27x <= 1204;
				I28x <= 1400;
				I29x <= 1540;
				I30x <= 1769;
				I31x <= 1916;
				I32x <= 2105;
				I33x <= 2285;
				I34x <= 2392;
				I35x <= 2433;
				I36x <= 2293;
				I37x <= 2015;
				I38x <= 1703;
				I39x <= 1368;
				I40x <= 1089;
				I41x <= 860;
				I42x <= 675;
				I43x <= 612;
				I44x <= 523;
				I45x <= 511;
				I46x <= 503;
				I47x <= 499;
				I48x <= 453;
				I49x <= 480;
				I50x <= 503;
				I51x <= 508;
				I52x <= 518;
				I53x <= 508;
				I54x <= 513;
				I55x <= 559;
				I56x <= 547;
				I57x <= 566;
				I58x <= 571;
				I59x <= 576;
				I60x <= 552;
				I61x <= 547;
				I62x <= 543;
				I63x <= 492;
				I64x <= 480;
				I65x <= 484;
				I66x <= 482;
				I67x <= 484;
				I68x <= 482;
				I69x <= 460;
				I70x <= 456;
				I71x <= 424;
				I72x <= 439;
				I73x <= 431;
				I74x <= 419;
				I75x <= 451;
				I76x <= 482;
				I77x <= 482;
				I78x <= 448;
				I79x <= 444;
				I80x <= 484;
				I81x <= 448;
				I82x <= 451;
				I83x <= 465;
				I84x <= 441;
				I85x <= 470;
				I86x <= 434;
				I87x <= 446;
				I88x <= 457;
				I89x <= 405;
				I90x <= 410;
				I91x <= 492;
				I92x <= 625;
				I93x <= 719;
				I94x <= 719;
				I95x <= 835;
				I96x <= 966;
				I97x <= 1007;
				I98x <= 1146;
				I99x <= 1048;
				I100x <= 958;
				I101x <= 757;
				I102x <= 499;
				I103x <= 335;
				I104x <= 313;
				I105x <= 284;
				I106x <= 272;
				I107x <= 245;
				I108x <= 267;
				I109x <= 234;
				I110x <= 250;
				I111x <= 248;
				I112x <= 140;
				I113x <= 0;
				I114x <= 1843;
				I115x <= 4694;
				I116x <= 7405;
				I117x <= 7372;
				I118x <= 1933;
				I119x <= 586;
				I120x <= 743;
				I121x <= 771;
				I122x <= 615;
				I123x <= 516;
				I124x <= 477;
				I125x <= 465;
				I126x <= 482;
				I127x <= 465;
				I128x <= 482;
				I129x <= 480;
				I130x <= 484;
				I131x <= 480;
				I132x <= 472;
				I133x <= 484;
				I134x <= 451;
				I135x <= 482;
				I136x <= 543;
				I137x <= 561;
				I138x <= 643;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101010:begin
				I0x <= 8159;
				I1x <= 4464;
				I2x <= 1990;
				I3x <= 182;
				I4x <= 0;
				I5x <= 1744;
				I6x <= 2031;
				I7x <= 2023;
				I8x <= 2383;
				I9x <= 2523;
				I10x <= 2539;
				I11x <= 2670;
				I12x <= 2629;
				I13x <= 2678;
				I14x <= 2842;
				I15x <= 2834;
				I16x <= 2891;
				I17x <= 3014;
				I18x <= 3063;
				I19x <= 3031;
				I20x <= 3153;
				I21x <= 3309;
				I22x <= 3448;
				I23x <= 3694;
				I24x <= 4055;
				I25x <= 4390;
				I26x <= 4710;
				I27x <= 4947;
				I28x <= 5120;
				I29x <= 5275;
				I30x <= 5316;
				I31x <= 5349;
				I32x <= 5054;
				I33x <= 4694;
				I34x <= 4235;
				I35x <= 3784;
				I36x <= 3391;
				I37x <= 3031;
				I38x <= 2777;
				I39x <= 2629;
				I40x <= 2539;
				I41x <= 2465;
				I42x <= 2596;
				I43x <= 2482;
				I44x <= 2482;
				I45x <= 2342;
				I46x <= 2383;
				I47x <= 2367;
				I48x <= 2375;
				I49x <= 2342;
				I50x <= 2416;
				I51x <= 2383;
				I52x <= 2564;
				I53x <= 2490;
				I54x <= 2367;
				I55x <= 2441;
				I56x <= 2498;
				I57x <= 2465;
				I58x <= 2473;
				I59x <= 2482;
				I60x <= 2416;
				I61x <= 2457;
				I62x <= 2334;
				I63x <= 2342;
				I64x <= 2392;
				I65x <= 2334;
				I66x <= 2326;
				I67x <= 2301;
				I68x <= 2277;
				I69x <= 2285;
				I70x <= 2203;
				I71x <= 2269;
				I72x <= 2260;
				I73x <= 2408;
				I74x <= 2318;
				I75x <= 2269;
				I76x <= 2293;
				I77x <= 2318;
				I78x <= 2277;
				I79x <= 2359;
				I80x <= 2269;
				I81x <= 2293;
				I82x <= 2351;
				I83x <= 2482;
				I84x <= 2686;
				I85x <= 3039;
				I86x <= 3088;
				I87x <= 3366;
				I88x <= 3612;
				I89x <= 3604;
				I90x <= 3538;
				I91x <= 3661;
				I92x <= 3276;
				I93x <= 2965;
				I94x <= 2654;
				I95x <= 2465;
				I96x <= 2351;
				I97x <= 2424;
				I98x <= 2351;
				I99x <= 2383;
				I100x <= 2383;
				I101x <= 2318;
				I102x <= 2416;
				I103x <= 2490;
				I104x <= 3555;
				I105x <= 3710;
				I106x <= 4677;
				I107x <= 7938;
				I108x <= 8192;
				I109x <= 3555;
				I110x <= 1777;
				I111x <= 51;
				I112x <= 697;
				I113x <= 2138;
				I114x <= 2408;
				I115x <= 2555;
				I116x <= 2752;
				I117x <= 2875;
				I118x <= 2940;
				I119x <= 3006;
				I120x <= 2965;
				I121x <= 3145;
				I122x <= 3178;
				I123x <= 3203;
				I124x <= 3276;
				I125x <= 3366;
				I126x <= 3514;
				I127x <= 3506;
				I128x <= 3670;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101011:begin
				I0x <= 8192;
				I1x <= 2457;
				I2x <= 80;
				I3x <= 2203;
				I4x <= 2039;
				I5x <= 2310;
				I6x <= 1810;
				I7x <= 1605;
				I8x <= 1531;
				I9x <= 1327;
				I10x <= 1155;
				I11x <= 1245;
				I12x <= 1753;
				I13x <= 1105;
				I14x <= 1318;
				I15x <= 843;
				I16x <= 1105;
				I17x <= 1327;
				I18x <= 1048;
				I19x <= 1179;
				I20x <= 1114;
				I21x <= 1245;
				I22x <= 1351;
				I23x <= 1228;
				I24x <= 1351;
				I25x <= 1769;
				I26x <= 2088;
				I27x <= 2318;
				I28x <= 2031;
				I29x <= 2244;
				I30x <= 2441;
				I31x <= 2859;
				I32x <= 2392;
				I33x <= 2711;
				I34x <= 2506;
				I35x <= 1777;
				I36x <= 1974;
				I37x <= 1351;
				I38x <= 1687;
				I39x <= 1146;
				I40x <= 1310;
				I41x <= 818;
				I42x <= 917;
				I43x <= 1015;
				I44x <= 1081;
				I45x <= 901;
				I46x <= 1048;
				I47x <= 843;
				I48x <= 1220;
				I49x <= 1089;
				I50x <= 692;
				I51x <= 1220;
				I52x <= 909;
				I53x <= 1794;
				I54x <= 1196;
				I55x <= 1179;
				I56x <= 1097;
				I57x <= 1155;
				I58x <= 1368;
				I59x <= 1146;
				I60x <= 1015;
				I61x <= 1400;
				I62x <= 1515;
				I63x <= 1220;
				I64x <= 1384;
				I65x <= 1228;
				I66x <= 1400;
				I67x <= 1843;
				I68x <= 2048;
				I69x <= 2220;
				I70x <= 2056;
				I71x <= 2523;
				I72x <= 2506;
				I73x <= 2121;
				I74x <= 1695;
				I75x <= 1376;
				I76x <= 991;
				I77x <= 925;
				I78x <= 757;
				I79x <= 892;
				I80x <= 389;
				I81x <= 1376;
				I82x <= 752;
				I83x <= 827;
				I84x <= 772;
				I85x <= 1245;
				I86x <= 0;
				I87x <= 2244;
				I88x <= 5988;
				I89x <= 5185;
				I90x <= 827;
				I91x <= 1179;
				I92x <= 1941;
				I93x <= 1613;
				I94x <= 1269;
				I95x <= 958;
				I96x <= 942;
				I97x <= 1351;
				I98x <= 1196;
				I99x <= 958;
				I100x <= 958;
				I101x <= 1384;
				I102x <= 1040;
				I103x <= 827;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101100:begin
				I0x <= 8118;
				I1x <= 4988;
				I2x <= 974;
				I3x <= 262;
				I4x <= 547;
				I5x <= 421;
				I6x <= 353;
				I7x <= 303;
				I8x <= 337;
				I9x <= 307;
				I10x <= 351;
				I11x <= 353;
				I12x <= 376;
				I13x <= 463;
				I14x <= 441;
				I15x <= 449;
				I16x <= 536;
				I17x <= 522;
				I18x <= 581;
				I19x <= 618;
				I20x <= 656;
				I21x <= 693;
				I22x <= 746;
				I23x <= 892;
				I24x <= 991;
				I25x <= 1081;
				I26x <= 1269;
				I27x <= 1359;
				I28x <= 1548;
				I29x <= 1736;
				I30x <= 1892;
				I31x <= 2088;
				I32x <= 2244;
				I33x <= 2367;
				I34x <= 2310;
				I35x <= 2113;
				I36x <= 1908;
				I37x <= 1548;
				I38x <= 1212;
				I39x <= 884;
				I40x <= 665;
				I41x <= 544;
				I42x <= 359;
				I43x <= 296;
				I44x <= 245;
				I45x <= 203;
				I46x <= 213;
				I47x <= 190;
				I48x <= 253;
				I49x <= 249;
				I50x <= 248;
				I51x <= 311;
				I52x <= 280;
				I53x <= 329;
				I54x <= 341;
				I55x <= 347;
				I56x <= 384;
				I57x <= 335;
				I58x <= 341;
				I59x <= 286;
				I60x <= 282;
				I61x <= 315;
				I62x <= 272;
				I63x <= 329;
				I64x <= 288;
				I65x <= 248;
				I66x <= 290;
				I67x <= 227;
				I68x <= 270;
				I69x <= 237;
				I70x <= 222;
				I71x <= 292;
				I72x <= 241;
				I73x <= 278;
				I74x <= 303;
				I75x <= 235;
				I76x <= 248;
				I77x <= 203;
				I78x <= 256;
				I79x <= 258;
				I80x <= 227;
				I81x <= 249;
				I82x <= 229;
				I83x <= 282;
				I84x <= 272;
				I85x <= 240;
				I86x <= 286;
				I87x <= 262;
				I88x <= 371;
				I89x <= 396;
				I90x <= 433;
				I91x <= 477;
				I92x <= 421;
				I93x <= 481;
				I94x <= 500;
				I95x <= 437;
				I96x <= 416;
				I97x <= 347;
				I98x <= 410;
				I99x <= 280;
				I100x <= 150;
				I101x <= 154;
				I102x <= 127;
				I103x <= 134;
				I104x <= 131;
				I105x <= 115;
				I106x <= 140;
				I107x <= 134;
				I108x <= 168;
				I109x <= 104;
				I110x <= 0;
				I111x <= 44;
				I112x <= 1613;
				I113x <= 4276;
				I114x <= 6602;
				I115x <= 8192;
				I116x <= 5300;
				I117x <= 1122;
				I118x <= 319;
				I119x <= 536;
				I120x <= 410;
				I121x <= 312;
				I122x <= 253;
				I123x <= 270;
				I124x <= 245;
				I125x <= 278;
				I126x <= 312;
				I127x <= 333;
				I128x <= 439;
				I129x <= 441;
				I130x <= 414;
				I131x <= 465;
				I132x <= 480;
				I133x <= 575;
				I134x <= 566;
				I135x <= 587;
				I136x <= 634;
				I137x <= 691;
				I138x <= 843;
				I139x <= 917;
				I140x <= 1040;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101101:begin
				I0x <= 8192;
				I1x <= 5865;
				I2x <= 3727;
				I3x <= 1957;
				I4x <= 1310;
				I5x <= 1548;
				I6x <= 1572;
				I7x <= 1564;
				I8x <= 1507;
				I9x <= 1466;
				I10x <= 1523;
				I11x <= 1531;
				I12x <= 1613;
				I13x <= 1622;
				I14x <= 1613;
				I15x <= 1679;
				I16x <= 1671;
				I17x <= 1744;
				I18x <= 1761;
				I19x <= 1802;
				I20x <= 1892;
				I21x <= 1933;
				I22x <= 2072;
				I23x <= 2146;
				I24x <= 2228;
				I25x <= 2392;
				I26x <= 2465;
				I27x <= 2621;
				I28x <= 2670;
				I29x <= 2719;
				I30x <= 2801;
				I31x <= 2793;
				I32x <= 2801;
				I33x <= 2654;
				I34x <= 2441;
				I35x <= 2252;
				I36x <= 2015;
				I37x <= 1884;
				I38x <= 1753;
				I39x <= 1638;
				I40x <= 1589;
				I41x <= 1523;
				I42x <= 1548;
				I43x <= 1531;
				I44x <= 1490;
				I45x <= 1531;
				I46x <= 1490;
				I47x <= 1531;
				I48x <= 1507;
				I49x <= 1499;
				I50x <= 1515;
				I51x <= 1499;
				I52x <= 1556;
				I53x <= 1556;
				I54x <= 1548;
				I55x <= 1556;
				I56x <= 1507;
				I57x <= 1548;
				I58x <= 1540;
				I59x <= 1507;
				I60x <= 1540;
				I61x <= 1474;
				I62x <= 1507;
				I63x <= 1482;
				I64x <= 1466;
				I65x <= 1482;
				I66x <= 1466;
				I67x <= 1507;
				I68x <= 1597;
				I69x <= 1646;
				I70x <= 1769;
				I71x <= 1712;
				I72x <= 1818;
				I73x <= 1908;
				I74x <= 1925;
				I75x <= 1925;
				I76x <= 1785;
				I77x <= 1605;
				I78x <= 1425;
				I79x <= 1351;
				I80x <= 1351;
				I81x <= 1277;
				I82x <= 1302;
				I83x <= 1294;
				I84x <= 1253;
				I85x <= 1269;
				I86x <= 1236;
				I87x <= 1310;
				I88x <= 1294;
				I89x <= 1196;
				I90x <= 338;
				I91x <= 0;
				I92x <= 1843;
				I93x <= 4554;
				I94x <= 7946;
				I95x <= 6283;
				I96x <= 3891;
				I97x <= 2220;
				I98x <= 1376;
				I99x <= 1540;
				I100x <= 1638;
				I101x <= 1572;
				I102x <= 1597;
				I103x <= 1556;
				I104x <= 1515;
				I105x <= 1564;
				I106x <= 1564;
				I107x <= 1613;
				I108x <= 1654;
				I109x <= 1671;
				I110x <= 1712;
				I111x <= 1736;
				I112x <= 1826;
				I113x <= 1835;
				I114x <= 1859;
				I115x <= 1949;
				I116x <= 2007;
				I117x <= 2146;
				I118x <= 2236;
				I119x <= 2334;
				I120x <= 2482;
				I121x <= 2572;
				I122x <= 2736;
				I123x <= 2777;
				I124x <= 2785;
				I125x <= 2842;
				I126x <= 2818;
				I127x <= 2760;
				I128x <= 2547;
				I129x <= 2326;
				I130x <= 2129;
				I131x <= 1933;
				I132x <= 1835;
				I133x <= 1712;
				I134x <= 1630;
				I135x <= 1613;
				I136x <= 1597;
				I137x <= 1605;
				I138x <= 1589;
				I139x <= 1572;
				I140x <= 1605;
				I141x <= 1589;
				I142x <= 1638;
				I143x <= 1622;
				I144x <= 1605;
				I145x <= 1605;
				I146x <= 1597;
				I147x <= 1630;
				I148x <= 1622;
				I149x <= 1589;
				I150x <= 1581;
				I151x <= 1581;
				I152x <= 1613;
				I153x <= 1572;
				I154x <= 1531;
				I155x <= 1548;
				I156x <= 1531;
				I157x <= 1581;
				I158x <= 1548;
				I159x <= 1507;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101110:begin
				I0x <= 7757;
				I1x <= 6717;
				I2x <= 3891;
				I3x <= 2031;
				I4x <= 1220;
				I5x <= 1474;
				I6x <= 1589;
				I7x <= 1523;
				I8x <= 1507;
				I9x <= 1572;
				I10x <= 1556;
				I11x <= 1589;
				I12x <= 1630;
				I13x <= 1622;
				I14x <= 1679;
				I15x <= 1720;
				I16x <= 1761;
				I17x <= 1794;
				I18x <= 1802;
				I19x <= 1875;
				I20x <= 1949;
				I21x <= 2048;
				I22x <= 2129;
				I23x <= 2236;
				I24x <= 2367;
				I25x <= 2523;
				I26x <= 2621;
				I27x <= 2752;
				I28x <= 2818;
				I29x <= 2859;
				I30x <= 2908;
				I31x <= 2891;
				I32x <= 2785;
				I33x <= 2605;
				I34x <= 2367;
				I35x <= 2129;
				I36x <= 1966;
				I37x <= 1851;
				I38x <= 1703;
				I39x <= 1613;
				I40x <= 1572;
				I41x <= 1548;
				I42x <= 1523;
				I43x <= 1523;
				I44x <= 1540;
				I45x <= 1490;
				I46x <= 1523;
				I47x <= 1515;
				I48x <= 1523;
				I49x <= 1564;
				I50x <= 1556;
				I51x <= 1540;
				I52x <= 1589;
				I53x <= 1597;
				I54x <= 1605;
				I55x <= 1622;
				I56x <= 1622;
				I57x <= 1613;
				I58x <= 1613;
				I59x <= 1613;
				I60x <= 1597;
				I61x <= 1548;
				I62x <= 1556;
				I63x <= 1548;
				I64x <= 1523;
				I65x <= 1523;
				I66x <= 1523;
				I67x <= 1523;
				I68x <= 1523;
				I69x <= 1482;
				I70x <= 1523;
				I71x <= 1654;
				I72x <= 1753;
				I73x <= 1826;
				I74x <= 1802;
				I75x <= 1867;
				I76x <= 1990;
				I77x <= 2015;
				I78x <= 2039;
				I79x <= 1925;
				I80x <= 1671;
				I81x <= 1482;
				I82x <= 1409;
				I83x <= 1368;
				I84x <= 1277;
				I85x <= 1261;
				I86x <= 1277;
				I87x <= 1269;
				I88x <= 1302;
				I89x <= 1286;
				I90x <= 1277;
				I91x <= 1294;
				I92x <= 1286;
				I93x <= 1089;
				I94x <= 0;
				I95x <= 116;
				I96x <= 2228;
				I97x <= 5259;
				I98x <= 8192;
				I99x <= 5865;
				I100x <= 3497;
				I101x <= 1646;
				I102x <= 1245;
				I103x <= 1507;
				I104x <= 1564;
				I105x <= 1523;
				I106x <= 1499;
				I107x <= 1523;
				I108x <= 1556;
				I109x <= 1564;
				I110x <= 1564;
				I111x <= 1597;
				I112x <= 1581;
				I113x <= 1630;
				I114x <= 1638;
				I115x <= 1703;
				I116x <= 1744;
				I117x <= 1802;
				I118x <= 1884;
				I119x <= 1990;
				I120x <= 2072;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00101111:begin
				I0x <= 8110;
				I1x <= 6447;
				I2x <= 3932;
				I3x <= 2170;
				I4x <= 1449;
				I5x <= 1728;
				I6x <= 1777;
				I7x <= 1712;
				I8x <= 1703;
				I9x <= 1728;
				I10x <= 1736;
				I11x <= 1769;
				I12x <= 1785;
				I13x <= 1794;
				I14x <= 1843;
				I15x <= 1851;
				I16x <= 1900;
				I17x <= 1933;
				I18x <= 1982;
				I19x <= 2039;
				I20x <= 2113;
				I21x <= 2179;
				I22x <= 2269;
				I23x <= 2383;
				I24x <= 2514;
				I25x <= 2670;
				I26x <= 2793;
				I27x <= 2916;
				I28x <= 3014;
				I29x <= 3072;
				I30x <= 3121;
				I31x <= 3162;
				I32x <= 3112;
				I33x <= 2957;
				I34x <= 2695;
				I35x <= 2441;
				I36x <= 2203;
				I37x <= 2031;
				I38x <= 1875;
				I39x <= 1777;
				I40x <= 1728;
				I41x <= 1679;
				I42x <= 1662;
				I43x <= 1671;
				I44x <= 1671;
				I45x <= 1638;
				I46x <= 1654;
				I47x <= 1662;
				I48x <= 1662;
				I49x <= 1662;
				I50x <= 1654;
				I51x <= 1654;
				I52x <= 1671;
				I53x <= 1662;
				I54x <= 1671;
				I55x <= 1671;
				I56x <= 1662;
				I57x <= 1671;
				I58x <= 1654;
				I59x <= 1662;
				I60x <= 1646;
				I61x <= 1630;
				I62x <= 1630;
				I63x <= 1613;
				I64x <= 1605;
				I65x <= 1605;
				I66x <= 1597;
				I67x <= 1564;
				I68x <= 1581;
				I69x <= 1572;
				I70x <= 1564;
				I71x <= 1548;
				I72x <= 1548;
				I73x <= 1540;
				I74x <= 1548;
				I75x <= 1679;
				I76x <= 1769;
				I77x <= 1835;
				I78x <= 1810;
				I79x <= 1900;
				I80x <= 2007;
				I81x <= 1990;
				I82x <= 2064;
				I83x <= 1941;
				I84x <= 1728;
				I85x <= 1499;
				I86x <= 1441;
				I87x <= 1392;
				I88x <= 1359;
				I89x <= 1327;
				I90x <= 1318;
				I91x <= 1318;
				I92x <= 1310;
				I93x <= 1294;
				I94x <= 1327;
				I95x <= 1318;
				I96x <= 1310;
				I97x <= 1179;
				I98x <= 181;
				I99x <= 0;
				I100x <= 2072;
				I101x <= 5029;
				I102x <= 8192;
				I103x <= 6135;
				I104x <= 3645;
				I105x <= 1851;
				I106x <= 1335;
				I107x <= 1581;
				I108x <= 1597;
				I109x <= 1548;
				I110x <= 1548;
				I111x <= 1556;
				I112x <= 1564;
				I113x <= 1572;
				I114x <= 1630;
				I115x <= 1630;
				I116x <= 1654;
				I117x <= 1695;
				I118x <= 1728;
				I119x <= 1761;
				I120x <= 1818;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110000:begin
				I0x <= 8192;
				I1x <= 7757;
				I2x <= 3170;
				I3x <= 711;
				I4x <= 724;
				I5x <= 1032;
				I6x <= 815;
				I7x <= 709;
				I8x <= 680;
				I9x <= 670;
				I10x <= 680;
				I11x <= 712;
				I12x <= 711;
				I13x <= 722;
				I14x <= 758;
				I15x <= 815;
				I16x <= 819;
				I17x <= 843;
				I18x <= 868;
				I19x <= 884;
				I20x <= 925;
				I21x <= 999;
				I22x <= 1024;
				I23x <= 1073;
				I24x <= 1163;
				I25x <= 1228;
				I26x <= 1327;
				I27x <= 1425;
				I28x <= 1556;
				I29x <= 1679;
				I30x <= 1785;
				I31x <= 1949;
				I32x <= 2072;
				I33x <= 2211;
				I34x <= 2301;
				I35x <= 2318;
				I36x <= 2252;
				I37x <= 2072;
				I38x <= 1843;
				I39x <= 1540;
				I40x <= 1318;
				I41x <= 1114;
				I42x <= 933;
				I43x <= 851;
				I44x <= 745;
				I45x <= 732;
				I46x <= 712;
				I47x <= 688;
				I48x <= 688;
				I49x <= 672;
				I50x <= 669;
				I51x <= 693;
				I52x <= 652;
				I53x <= 663;
				I54x <= 666;
				I55x <= 669;
				I56x <= 684;
				I57x <= 663;
				I58x <= 672;
				I59x <= 680;
				I60x <= 653;
				I61x <= 686;
				I62x <= 642;
				I63x <= 647;
				I64x <= 620;
				I65x <= 636;
				I66x <= 647;
				I67x <= 603;
				I68x <= 620;
				I69x <= 598;
				I70x <= 594;
				I71x <= 594;
				I72x <= 577;
				I73x <= 580;
				I74x <= 577;
				I75x <= 567;
				I76x <= 552;
				I77x <= 533;
				I78x <= 546;
				I79x <= 523;
				I80x <= 539;
				I81x <= 537;
				I82x <= 497;
				I83x <= 544;
				I84x <= 523;
				I85x <= 525;
				I86x <= 529;
				I87x <= 525;
				I88x <= 550;
				I89x <= 531;
				I90x <= 516;
				I91x <= 529;
				I92x <= 520;
				I93x <= 533;
				I94x <= 531;
				I95x <= 493;
				I96x <= 514;
				I97x <= 485;
				I98x <= 508;
				I99x <= 500;
				I100x <= 483;
				I101x <= 512;
				I102x <= 474;
				I103x <= 516;
				I104x <= 468;
				I105x <= 485;
				I106x <= 523;
				I107x <= 453;
				I108x <= 497;
				I109x <= 480;
				I110x <= 483;
				I111x <= 500;
				I112x <= 523;
				I113x <= 625;
				I114x <= 676;
				I115x <= 892;
				I116x <= 942;
				I117x <= 901;
				I118x <= 1081;
				I119x <= 1073;
				I120x <= 1007;
				I121x <= 950;
				I122x <= 791;
				I123x <= 675;
				I124x <= 602;
				I125x <= 448;
				I126x <= 424;
				I127x <= 389;
				I128x <= 401;
				I129x <= 353;
				I130x <= 371;
				I131x <= 378;
				I132x <= 374;
				I133x <= 97;
				I134x <= 0;
				I135x <= 810;
				I136x <= 3334;
				I137x <= 7487;
				I138x <= 8118;
				I139x <= 3842;
				I140x <= 892;
				I141x <= 603;
				I142x <= 843;
				I143x <= 680;
				I144x <= 577;
				I145x <= 546;
				I146x <= 543;
				I147x <= 577;
				I148x <= 579;
				I149x <= 590;
				I150x <= 630;
				I151x <= 655;
				I152x <= 636;
				I153x <= 699;
				I154x <= 726;
				I155x <= 747;
				I156x <= 792;
				I157x <= 804;
				I158x <= 884;
				I159x <= 892;
				I160x <= 974;
				I161x <= 1048;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110001:begin
				I0x <= 7389;
				I1x <= 8192;
				I2x <= 3055;
				I3x <= 1122;
				I4x <= 1048;
				I5x <= 860;
				I6x <= 925;
				I7x <= 851;
				I8x <= 835;
				I9x <= 860;
				I10x <= 851;
				I11x <= 835;
				I12x <= 790;
				I13x <= 813;
				I14x <= 868;
				I15x <= 884;
				I16x <= 933;
				I17x <= 917;
				I18x <= 999;
				I19x <= 1105;
				I20x <= 1212;
				I21x <= 1318;
				I22x <= 1425;
				I23x <= 1622;
				I24x <= 1867;
				I25x <= 2105;
				I26x <= 2375;
				I27x <= 2596;
				I28x <= 2826;
				I29x <= 3014;
				I30x <= 3162;
				I31x <= 3268;
				I32x <= 3137;
				I33x <= 2916;
				I34x <= 2572;
				I35x <= 2228;
				I36x <= 1835;
				I37x <= 1515;
				I38x <= 1253;
				I39x <= 1056;
				I40x <= 966;
				I41x <= 851;
				I42x <= 779;
				I43x <= 770;
				I44x <= 770;
				I45x <= 763;
				I46x <= 705;
				I47x <= 759;
				I48x <= 763;
				I49x <= 724;
				I50x <= 736;
				I51x <= 736;
				I52x <= 716;
				I53x <= 736;
				I54x <= 651;
				I55x <= 666;
				I56x <= 628;
				I57x <= 585;
				I58x <= 589;
				I59x <= 520;
				I60x <= 551;
				I61x <= 478;
				I62x <= 501;
				I63x <= 501;
				I64x <= 393;
				I65x <= 493;
				I66x <= 431;
				I67x <= 385;
				I68x <= 389;
				I69x <= 416;
				I70x <= 443;
				I71x <= 412;
				I72x <= 358;
				I73x <= 358;
				I74x <= 331;
				I75x <= 320;
				I76x <= 335;
				I77x <= 254;
				I78x <= 312;
				I79x <= 300;
				I80x <= 339;
				I81x <= 331;
				I82x <= 308;
				I83x <= 373;
				I84x <= 366;
				I85x <= 512;
				I86x <= 675;
				I87x <= 736;
				I88x <= 843;
				I89x <= 1048;
				I90x <= 999;
				I91x <= 868;
				I92x <= 797;
				I93x <= 728;
				I94x <= 420;
				I95x <= 408;
				I96x <= 192;
				I97x <= 150;
				I98x <= 235;
				I99x <= 227;
				I100x <= 0;
				I101x <= 123;
				I102x <= 2154;
				I103x <= 5103;
				I104x <= 6881;
				I105x <= 6094;
				I106x <= 1417;
				I107x <= 659;
				I108x <= 381;
				I109x <= 335;
				I110x <= 389;
				I111x <= 273;
				I112x <= 304;
				I113x <= 277;
				I114x <= 281;
				I115x <= 331;
				I116x <= 242;
				I117x <= 293;
				I118x <= 354;
				I119x <= 343;
				I120x <= 370;
				I121x <= 420;
				I122x <= 443;
				I123x <= 574;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110010:begin
				I0x <= 8132;
				I1x <= 8109;
				I2x <= 5307;
				I3x <= 4138;
				I4x <= 3299;
				I5x <= 2866;
				I6x <= 2242;
				I7x <= 2027;
				I8x <= 1750;
				I9x <= 1717;
				I10x <= 1714;
				I11x <= 1694;
				I12x <= 1642;
				I13x <= 1615;
				I14x <= 1719;
				I15x <= 1687;
				I16x <= 1638;
				I17x <= 1629;
				I18x <= 1579;
				I19x <= 1541;
				I20x <= 1482;
				I21x <= 1442;
				I22x <= 1458;
				I23x <= 1424;
				I24x <= 1383;
				I25x <= 1343;
				I26x <= 1300;
				I27x <= 1345;
				I28x <= 1357;
				I29x <= 1370;
				I30x <= 1485;
				I31x <= 1482;
				I32x <= 1615;
				I33x <= 1752;
				I34x <= 1883;
				I35x <= 1953;
				I36x <= 2072;
				I37x <= 2157;
				I38x <= 2198;
				I39x <= 2184;
				I40x <= 2137;
				I41x <= 2123;
				I42x <= 2094;
				I43x <= 2121;
				I44x <= 2016;
				I45x <= 1957;
				I46x <= 1937;
				I47x <= 1923;
				I48x <= 1867;
				I49x <= 1826;
				I50x <= 1878;
				I51x <= 1818;
				I52x <= 1826;
				I53x <= 1854;
				I54x <= 1815;
				I55x <= 1835;
				I56x <= 1804;
				I57x <= 1766;
				I58x <= 1844;
				I59x <= 1835;
				I60x <= 1905;
				I61x <= 1912;
				I62x <= 1903;
				I63x <= 2007;
				I64x <= 2029;
				I65x <= 1979;
				I66x <= 1998;
				I67x <= 1975;
				I68x <= 1883;
				I69x <= 1959;
				I70x <= 1881;
				I71x <= 1943;
				I72x <= 1953;
				I73x <= 1970;
				I74x <= 1939;
				I75x <= 2043;
				I76x <= 2033;
				I77x <= 1988;
				I78x <= 2263;
				I79x <= 2342;
				I80x <= 2170;
				I81x <= 2227;
				I82x <= 2202;
				I83x <= 2087;
				I84x <= 1831;
				I85x <= 1806;
				I86x <= 1788;
				I87x <= 1849;
				I88x <= 1800;
				I89x <= 1876;
				I90x <= 1876;
				I91x <= 1862;
				I92x <= 1437;
				I93x <= 477;
				I94x <= 0;
				I95x <= 551;
				I96x <= 1489;
				I97x <= 2942;
				I98x <= 4496;
				I99x <= 5624;
				I100x <= 7621;
				I101x <= 8192;
				I102x <= 7388;
				I103x <= 4383;
				I104x <= 3324;
				I105x <= 2712;
				I106x <= 2411;
				I107x <= 2083;
				I108x <= 2045;
				I109x <= 2043;
				I110x <= 2015;
				I111x <= 1959;
				I112x <= 1973;
				I113x <= 1957;
				I114x <= 1919;
				I115x <= 1899;
				I116x <= 1865;
				I117x <= 1860;
				I118x <= 1815;
				I119x <= 1775;
				I120x <= 1730;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110011:begin
				I0x <= 8192;
				I1x <= 7131;
				I2x <= 5566;
				I3x <= 3322;
				I4x <= 186;
				I5x <= 363;
				I6x <= 745;
				I7x <= 1357;
				I8x <= 1490;
				I9x <= 1441;
				I10x <= 1561;
				I11x <= 1383;
				I12x <= 1698;
				I13x <= 1694;
				I14x <= 1534;
				I15x <= 1734;
				I16x <= 1516;
				I17x <= 1853;
				I18x <= 1849;
				I19x <= 1769;
				I20x <= 1982;
				I21x <= 1805;
				I22x <= 2102;
				I23x <= 2177;
				I24x <= 1885;
				I25x <= 2270;
				I26x <= 2040;
				I27x <= 2266;
				I28x <= 2368;
				I29x <= 2315;
				I30x <= 2616;
				I31x <= 2306;
				I32x <= 2550;
				I33x <= 2585;
				I34x <= 2434;
				I35x <= 2585;
				I36x <= 2262;
				I37x <= 2332;
				I38x <= 2222;
				I39x <= 1902;
				I40x <= 2000;
				I41x <= 1494;
				I42x <= 1760;
				I43x <= 1685;
				I44x <= 1463;
				I45x <= 1729;
				I46x <= 1405;
				I47x <= 1578;
				I48x <= 1707;
				I49x <= 1578;
				I50x <= 1747;
				I51x <= 1379;
				I52x <= 1680;
				I53x <= 1694;
				I54x <= 1539;
				I55x <= 1720;
				I56x <= 1463;
				I57x <= 1676;
				I58x <= 1636;
				I59x <= 1468;
				I60x <= 1725;
				I61x <= 1312;
				I62x <= 1618;
				I63x <= 1623;
				I64x <= 1472;
				I65x <= 1556;
				I66x <= 1250;
				I67x <= 1508;
				I68x <= 1530;
				I69x <= 1321;
				I70x <= 1516;
				I71x <= 1131;
				I72x <= 1370;
				I73x <= 1374;
				I74x <= 1193;
				I75x <= 1339;
				I76x <= 1117;
				I77x <= 1352;
				I78x <= 1303;
				I79x <= 1179;
				I80x <= 1423;
				I81x <= 1188;
				I82x <= 1561;
				I83x <= 1751;
				I84x <= 1623;
				I85x <= 1836;
				I86x <= 1902;
				I87x <= 2364;
				I88x <= 2208;
				I89x <= 2066;
				I90x <= 1765;
				I91x <= 1317;
				I92x <= 1423;
				I93x <= 1122;
				I94x <= 820;
				I95x <= 873;
				I96x <= 669;
				I97x <= 860;
				I98x <= 820;
				I99x <= 687;
				I100x <= 824;
				I101x <= 0;
				I102x <= 1028;
				I103x <= 2807;
				I104x <= 5109;
				I105x <= 7770;
				I106x <= 7726;
				I107x <= 5619;
				I108x <= 3534;
				I109x <= 359;
				I110x <= 221;
				I111x <= 660;
				I112x <= 1095;
				I113x <= 1264;
				I114x <= 1268;
				I115x <= 1521;
				I116x <= 1241;
				I117x <= 1476;
				I118x <= 1459;
				I119x <= 1397;
				I120x <= 1663;
				I121x <= 1330;
				I122x <= 1601;
				I123x <= 1578;
				I124x <= 1556;
				I125x <= 1809;
				I126x <= 1556;
				I127x <= 1889;
				I128x <= 1849;
				I129x <= 1787;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110100:begin
				I0x <= 8123;
				I1x <= 6476;
				I2x <= 1974;
				I3x <= 1479;
				I4x <= 1103;
				I5x <= 901;
				I6x <= 778;
				I7x <= 689;
				I8x <= 785;
				I9x <= 727;
				I10x <= 707;
				I11x <= 698;
				I12x <= 680;
				I13x <= 678;
				I14x <= 707;
				I15x <= 729;
				I16x <= 685;
				I17x <= 680;
				I18x <= 687;
				I19x <= 616;
				I20x <= 816;
				I21x <= 887;
				I22x <= 914;
				I23x <= 1043;
				I24x <= 1057;
				I25x <= 1132;
				I26x <= 1304;
				I27x <= 1290;
				I28x <= 1466;
				I29x <= 1568;
				I30x <= 1722;
				I31x <= 1945;
				I32x <= 1811;
				I33x <= 1911;
				I34x <= 1956;
				I35x <= 2089;
				I36x <= 1976;
				I37x <= 1675;
				I38x <= 1546;
				I39x <= 1297;
				I40x <= 1099;
				I41x <= 950;
				I42x <= 843;
				I43x <= 761;
				I44x <= 734;
				I45x <= 674;
				I46x <= 689;
				I47x <= 707;
				I48x <= 736;
				I49x <= 627;
				I50x <= 689;
				I51x <= 743;
				I52x <= 652;
				I53x <= 816;
				I54x <= 749;
				I55x <= 821;
				I56x <= 796;
				I57x <= 761;
				I58x <= 876;
				I59x <= 770;
				I60x <= 794;
				I61x <= 763;
				I62x <= 680;
				I63x <= 792;
				I64x <= 765;
				I65x <= 756;
				I66x <= 596;
				I67x <= 752;
				I68x <= 734;
				I69x <= 810;
				I70x <= 734;
				I71x <= 685;
				I72x <= 741;
				I73x <= 732;
				I74x <= 689;
				I75x <= 658;
				I76x <= 680;
				I77x <= 685;
				I78x <= 645;
				I79x <= 770;
				I80x <= 879;
				I81x <= 968;
				I82x <= 934;
				I83x <= 870;
				I84x <= 787;
				I85x <= 638;
				I86x <= 736;
				I87x <= 758;
				I88x <= 747;
				I89x <= 603;
				I90x <= 449;
				I91x <= 413;
				I92x <= 433;
				I93x <= 362;
				I94x <= 358;
				I95x <= 505;
				I96x <= 478;
				I97x <= 0;
				I98x <= 1404;
				I99x <= 3382;
				I100x <= 6062;
				I101x <= 7680;
				I102x <= 8192;
				I103x <= 4642;
				I104x <= 1439;
				I105x <= 1163;
				I106x <= 959;
				I107x <= 709;
				I108x <= 574;
				I109x <= 545;
				I110x <= 587;
				I111x <= 485;
				I112x <= 511;
				I113x <= 485;
				I114x <= 496;
				I115x <= 571;
				I116x <= 674;
				I117x <= 636;
				I118x <= 707;
				I119x <= 718;
				I120x <= 663;
				I121x <= 747;
				I122x <= 716;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110101:begin
				I0x <= 8192;
				I1x <= 6186;
				I2x <= 1582;
				I3x <= 0;
				I4x <= 1041;
				I5x <= 609;
				I6x <= 609;
				I7x <= 682;
				I8x <= 818;
				I9x <= 1123;
				I10x <= 937;
				I11x <= 1078;
				I12x <= 1050;
				I13x <= 1005;
				I14x <= 1219;
				I15x <= 1091;
				I16x <= 1191;
				I17x <= 1182;
				I18x <= 1109;
				I19x <= 1419;
				I20x <= 1237;
				I21x <= 1405;
				I22x <= 1441;
				I23x <= 1373;
				I24x <= 1651;
				I25x <= 1546;
				I26x <= 1687;
				I27x <= 1837;
				I28x <= 1805;
				I29x <= 2133;
				I30x <= 1992;
				I31x <= 2128;
				I32x <= 2196;
				I33x <= 2078;
				I34x <= 2278;
				I35x <= 2110;
				I36x <= 2119;
				I37x <= 2042;
				I38x <= 1814;
				I39x <= 1992;
				I40x <= 1728;
				I41x <= 1783;
				I42x <= 1746;
				I43x <= 1582;
				I44x <= 1746;
				I45x <= 1587;
				I46x <= 1673;
				I47x <= 1569;
				I48x <= 1441;
				I49x <= 1669;
				I50x <= 1532;
				I51x <= 1601;
				I52x <= 1505;
				I53x <= 1355;
				I54x <= 1610;
				I55x <= 1414;
				I56x <= 1464;
				I57x <= 1432;
				I58x <= 1282;
				I59x <= 1541;
				I60x <= 1391;
				I61x <= 1473;
				I62x <= 1460;
				I63x <= 1314;
				I64x <= 1491;
				I65x <= 1464;
				I66x <= 1537;
				I67x <= 1528;
				I68x <= 1491;
				I69x <= 1792;
				I70x <= 1664;
				I71x <= 1760;
				I72x <= 1696;
				I73x <= 1610;
				I74x <= 1664;
				I75x <= 1246;
				I76x <= 987;
				I77x <= 1237;
				I78x <= 1064;
				I79x <= 1541;
				I80x <= 1259;
				I81x <= 1187;
				I82x <= 1168;
				I83x <= 1364;
				I84x <= 2983;
				I85x <= 4189;
				I86x <= 5058;
				I87x <= 7063;
				I88x <= 7832;
				I89x <= 3939;
				I90x <= 450;
				I91x <= 90;
				I92x <= 632;
				I93x <= 450;
				I94x <= 809;
				I95x <= 727;
				I96x <= 877;
				I97x <= 864;
				I98x <= 755;
				I99x <= 1114;
				I100x <= 1023;
				I101x <= 1059;
				I102x <= 1005;
				I103x <= 882;
				I104x <= 1246;
				I105x <= 1141;
				I106x <= 1219;
				I107x <= 1173;
				I108x <= 1041;
				I109x <= 1428;
				I110x <= 1350;
				I111x <= 1432;
				I112x <= 1473;
				I113x <= 1341;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110110:begin
				I0x <= 8192;
				I1x <= 5237;
				I2x <= 2547;
				I3x <= 1017;
				I4x <= 152;
				I5x <= 666;
				I6x <= 701;
				I7x <= 915;
				I8x <= 935;
				I9x <= 706;
				I10x <= 935;
				I11x <= 894;
				I12x <= 996;
				I13x <= 1139;
				I14x <= 747;
				I15x <= 1174;
				I16x <= 1067;
				I17x <= 1052;
				I18x <= 991;
				I19x <= 874;
				I20x <= 1017;
				I21x <= 1108;
				I22x <= 1062;
				I23x <= 1235;
				I24x <= 1108;
				I25x <= 1357;
				I26x <= 1133;
				I27x <= 1469;
				I28x <= 1383;
				I29x <= 1220;
				I30x <= 1301;
				I31x <= 1398;
				I32x <= 1184;
				I33x <= 1245;
				I34x <= 762;
				I35x <= 823;
				I36x <= 594;
				I37x <= 371;
				I38x <= 477;
				I39x <= 0;
				I40x <= 325;
				I41x <= 254;
				I42x <= 335;
				I43x <= 605;
				I44x <= 376;
				I45x <= 722;
				I46x <= 874;
				I47x <= 1011;
				I48x <= 1164;
				I49x <= 1001;
				I50x <= 1286;
				I51x <= 1286;
				I52x <= 1332;
				I53x <= 1515;
				I54x <= 1383;
				I55x <= 1576;
				I56x <= 1566;
				I57x <= 1428;
				I58x <= 1586;
				I59x <= 1388;
				I60x <= 1505;
				I61x <= 1540;
				I62x <= 1291;
				I63x <= 1617;
				I64x <= 1235;
				I65x <= 1398;
				I66x <= 1576;
				I67x <= 1454;
				I68x <= 1525;
				I69x <= 1220;
				I70x <= 1398;
				I71x <= 1306;
				I72x <= 1408;
				I73x <= 1495;
				I74x <= 1093;
				I75x <= 1357;
				I76x <= 1423;
				I77x <= 1439;
				I78x <= 1525;
				I79x <= 1342;
				I80x <= 1393;
				I81x <= 1210;
				I82x <= 1413;
				I83x <= 1464;
				I84x <= 1118;
				I85x <= 1449;
				I86x <= 1281;
				I87x <= 1378;
				I88x <= 1469;
				I89x <= 1276;
				I90x <= 1505;
				I91x <= 1744;
				I92x <= 2028;
				I93x <= 2120;
				I94x <= 2583;
				I95x <= 2878;
				I96x <= 2751;
				I97x <= 2959;
				I98x <= 3030;
				I99x <= 2303;
				I100x <= 1871;
				I101x <= 1561;
				I102x <= 1352;
				I103x <= 1296;
				I104x <= 1072;
				I105x <= 1281;
				I106x <= 1357;
				I107x <= 1210;
				I108x <= 1383;
				I109x <= 1047;
				I110x <= 711;
				I111x <= 1281;
				I112x <= 2257;
				I113x <= 5857;
				I114x <= 8136;
				I115x <= 4612;
				I116x <= 2918;
				I117x <= 1550;
				I118x <= 1205;
				I119x <= 1337;
				I120x <= 1576;
				I121x <= 1586;
				I122x <= 1571;
				I123x <= 1601;
				I124x <= 1342;
				I125x <= 1667;
				I126x <= 1632;
				I127x <= 1678;
				I128x <= 1800;
				I129x <= 1484;
				I130x <= 1779;
				I131x <= 1850;
				I132x <= 1784;
				I133x <= 1922;
				I134x <= 1688;
				I135x <= 1825;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00110111:begin
				I0x <= 7825;
				I1x <= 6835;
				I2x <= 4011;
				I3x <= 3814;
				I4x <= 3488;
				I5x <= 2805;
				I6x <= 3007;
				I7x <= 3076;
				I8x <= 2764;
				I9x <= 2768;
				I10x <= 3043;
				I11x <= 2929;
				I12x <= 3062;
				I13x <= 3364;
				I14x <= 3341;
				I15x <= 3268;
				I16x <= 3025;
				I17x <= 3227;
				I18x <= 3314;
				I19x <= 3259;
				I20x <= 3451;
				I21x <= 3603;
				I22x <= 3484;
				I23x <= 3250;
				I24x <= 3571;
				I25x <= 3410;
				I26x <= 3383;
				I27x <= 3474;
				I28x <= 3318;
				I29x <= 3511;
				I30x <= 2929;
				I31x <= 3181;
				I32x <= 2970;
				I33x <= 3021;
				I34x <= 2952;
				I35x <= 2608;
				I36x <= 2782;
				I37x <= 3108;
				I38x <= 2668;
				I39x <= 2736;
				I40x <= 2819;
				I41x <= 3007;
				I42x <= 2727;
				I43x <= 3025;
				I44x <= 2571;
				I45x <= 2723;
				I46x <= 2791;
				I47x <= 2686;
				I48x <= 2842;
				I49x <= 2732;
				I50x <= 2700;
				I51x <= 2791;
				I52x <= 2415;
				I53x <= 2814;
				I54x <= 2443;
				I55x <= 2470;
				I56x <= 2489;
				I57x <= 2493;
				I58x <= 2956;
				I59x <= 2709;
				I60x <= 2535;
				I61x <= 2883;
				I62x <= 3043;
				I63x <= 3218;
				I64x <= 3479;
				I65x <= 3539;
				I66x <= 4002;
				I67x <= 3901;
				I68x <= 3965;
				I69x <= 3699;
				I70x <= 3479;
				I71x <= 3163;
				I72x <= 2865;
				I73x <= 2191;
				I74x <= 2521;
				I75x <= 2205;
				I76x <= 2447;
				I77x <= 2260;
				I78x <= 1618;
				I79x <= 265;
				I80x <= 0;
				I81x <= 3804;
				I82x <= 7146;
				I83x <= 8192;
				I84x <= 6917;
				I85x <= 4098;
				I86x <= 3575;
				I87x <= 2622;
				I88x <= 3263;
				I89x <= 3158;
				I90x <= 2755;
				I91x <= 2768;
				I92x <= 2910;
				I93x <= 2764;
				I94x <= 2933;
				I95x <= 2938;
				I96x <= 3231;
				I97x <= 3131;
				I98x <= 3094;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111000:begin
				I0x <= 8168;
				I1x <= 8192;
				I2x <= 8105;
				I3x <= 7728;
				I4x <= 7246;
				I5x <= 6812;
				I6x <= 6301;
				I7x <= 6000;
				I8x <= 5542;
				I9x <= 5055;
				I10x <= 5038;
				I11x <= 4852;
				I12x <= 4725;
				I13x <= 4812;
				I14x <= 4962;
				I15x <= 4823;
				I16x <= 4922;
				I17x <= 4748;
				I18x <= 4742;
				I19x <= 4829;
				I20x <= 4754;
				I21x <= 4730;
				I22x <= 4701;
				I23x <= 4632;
				I24x <= 4638;
				I25x <= 4638;
				I26x <= 4446;
				I27x <= 4382;
				I28x <= 4487;
				I29x <= 4516;
				I30x <= 4504;
				I31x <= 4377;
				I32x <= 4330;
				I33x <= 4330;
				I34x <= 4330;
				I35x <= 4336;
				I36x <= 4261;
				I37x <= 4156;
				I38x <= 4371;
				I39x <= 4191;
				I40x <= 4435;
				I41x <= 4516;
				I42x <= 4591;
				I43x <= 4840;
				I44x <= 4742;
				I45x <= 4777;
				I46x <= 5443;
				I47x <= 5345;
				I48x <= 5559;
				I49x <= 5704;
				I50x <= 5646;
				I51x <= 5432;
				I52x <= 4887;
				I53x <= 4440;
				I54x <= 4133;
				I55x <= 3866;
				I56x <= 3832;
				I57x <= 3577;
				I58x <= 3455;
				I59x <= 3495;
				I60x <= 3351;
				I61x <= 3490;
				I62x <= 3530;
				I63x <= 3809;
				I64x <= 4185;
				I65x <= 4632;
				I66x <= 6806;
				I67x <= 7136;
				I68x <= 3513;
				I69x <= 0;
				I70x <= 626;
				I71x <= 1750;
				I72x <= 2533;
				I73x <= 3223;
				I74x <= 3449;
				I75x <= 3710;
				I76x <= 3791;
				I77x <= 3693;
				I78x <= 3774;
				I79x <= 3774;
				I80x <= 3849;
				I81x <= 3710;
				I82x <= 3924;
				I83x <= 4098;
				I84x <= 4156;
				I85x <= 4249;
				I86x <= 4435;
				I87x <= 4452;
				I88x <= 4614;
				I89x <= 4887;
				I90x <= 4997;
				I91x <= 5385;
				I92x <= 5722;
				I93x <= 6029;
				I94x <= 6452;
				I95x <= 6806;
				I96x <= 7044;
				I97x <= 7490;
				I98x <= 7525;
				I99x <= 7670;
				I100x <= 7583;
				I101x <= 7531;
				I102x <= 7333;
				I103x <= 6858;
				I104x <= 6435;
				I105x <= 5872;
				I106x <= 5693;
				I107x <= 5252;
				I108x <= 4893;
				I109x <= 4806;
				I110x <= 4574;
				I111x <= 4522;
				I112x <= 4527;
				I113x <= 4667;
				I114x <= 4475;
				I115x <= 4464;
				I116x <= 4545;
				I117x <= 4440;
				I118x <= 4527;
				I119x <= 4342;
				I120x <= 4359;
				I121x <= 4382;
				I122x <= 4069;
				I123x <= 4278;
				I124x <= 4267;
				I125x <= 4336;
				I126x <= 4284;
				I127x <= 4353;
				I128x <= 4411;
				I129x <= 4417;
				I130x <= 4209;
				I131x <= 4238;
				I132x <= 4336;
				I133x <= 4313;
				I134x <= 4243;
				I135x <= 4220;
				I136x <= 4046;
				I137x <= 4023;
				I138x <= 4180;
				I139x <= 4353;
				I140x <= 4562;
				I141x <= 4655;
				I142x <= 4690;
				I143x <= 4875;
				I144x <= 4881;
				I145x <= 5142;
				I146x <= 5432;
				I147x <= 5345;
				I148x <= 5791;
				I149x <= 5333;
				I150x <= 5757;
				I151x <= 5183;
				I152x <= 4684;
				I153x <= 4446;
				I154x <= 4191;
				I155x <= 4104;
				I156x <= 3872;
				I157x <= 3646;
				I158x <= 3727;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111001:begin
				I0x <= 7978;
				I1x <= 5437;
				I2x <= 2804;
				I3x <= 1393;
				I4x <= 1368;
				I5x <= 2214;
				I6x <= 2913;
				I7x <= 2708;
				I8x <= 2959;
				I9x <= 2838;
				I10x <= 2733;
				I11x <= 3034;
				I12x <= 3009;
				I13x <= 3114;
				I14x <= 3202;
				I15x <= 3097;
				I16x <= 3202;
				I17x <= 3160;
				I18x <= 3193;
				I19x <= 3135;
				I20x <= 3219;
				I21x <= 3491;
				I22x <= 3235;
				I23x <= 3415;
				I24x <= 3411;
				I25x <= 3570;
				I26x <= 3834;
				I27x <= 3796;
				I28x <= 3809;
				I29x <= 3851;
				I30x <= 3846;
				I31x <= 3779;
				I32x <= 3759;
				I33x <= 3796;
				I34x <= 3495;
				I35x <= 3252;
				I36x <= 3256;
				I37x <= 3047;
				I38x <= 2821;
				I39x <= 2842;
				I40x <= 2704;
				I41x <= 2653;
				I42x <= 2796;
				I43x <= 2741;
				I44x <= 2632;
				I45x <= 2553;
				I46x <= 2896;
				I47x <= 2766;
				I48x <= 2833;
				I49x <= 2653;
				I50x <= 2699;
				I51x <= 2624;
				I52x <= 2729;
				I53x <= 2733;
				I54x <= 2528;
				I55x <= 2503;
				I56x <= 2666;
				I57x <= 2515;
				I58x <= 2519;
				I59x <= 2423;
				I60x <= 2507;
				I61x <= 2545;
				I62x <= 2411;
				I63x <= 2683;
				I64x <= 2511;
				I65x <= 2319;
				I66x <= 2310;
				I67x <= 2486;
				I68x <= 2708;
				I69x <= 2829;
				I70x <= 2829;
				I71x <= 2892;
				I72x <= 2787;
				I73x <= 3051;
				I74x <= 2867;
				I75x <= 2490;
				I76x <= 2666;
				I77x <= 2406;
				I78x <= 2499;
				I79x <= 2231;
				I80x <= 2235;
				I81x <= 2113;
				I82x <= 2201;
				I83x <= 2026;
				I84x <= 581;
				I85x <= 0;
				I86x <= 1213;
				I87x <= 4545;
				I88x <= 8192;
				I89x <= 6630;
				I90x <= 3101;
				I91x <= 1557;
				I92x <= 1486;
				I93x <= 2285;
				I94x <= 2482;
				I95x <= 2632;
				I96x <= 2783;
				I97x <= 2729;
				I98x <= 2771;
				I99x <= 2716;
				I100x <= 2938;
				I101x <= 3005;
				I102x <= 2892;
				I103x <= 2959;
				I104x <= 3030;
				I105x <= 3034;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111010:begin
				I0x <= 7909;
				I1x <= 3966;
				I2x <= 778;
				I3x <= 173;
				I4x <= 0;
				I5x <= 459;
				I6x <= 695;
				I7x <= 891;
				I8x <= 931;
				I9x <= 968;
				I10x <= 1084;
				I11x <= 1064;
				I12x <= 1117;
				I13x <= 1181;
				I14x <= 1307;
				I15x <= 1314;
				I16x <= 1337;
				I17x <= 1374;
				I18x <= 1487;
				I19x <= 1630;
				I20x <= 1693;
				I21x <= 1716;
				I22x <= 1820;
				I23x <= 2122;
				I24x <= 2136;
				I25x <= 2239;
				I26x <= 2222;
				I27x <= 2352;
				I28x <= 2299;
				I29x <= 2186;
				I30x <= 1933;
				I31x <= 1800;
				I32x <= 1700;
				I33x <= 1686;
				I34x <= 1310;
				I35x <= 1301;
				I36x <= 1221;
				I37x <= 1154;
				I38x <= 981;
				I39x <= 1044;
				I40x <= 1154;
				I41x <= 1151;
				I42x <= 1117;
				I43x <= 1224;
				I44x <= 1284;
				I45x <= 1384;
				I46x <= 1400;
				I47x <= 1400;
				I48x <= 1500;
				I49x <= 1261;
				I50x <= 1460;
				I51x <= 1487;
				I52x <= 1414;
				I53x <= 1493;
				I54x <= 1294;
				I55x <= 1370;
				I56x <= 1157;
				I57x <= 1211;
				I58x <= 1201;
				I59x <= 1161;
				I60x <= 1281;
				I61x <= 1424;
				I62x <= 1587;
				I63x <= 1753;
				I64x <= 1733;
				I65x <= 1743;
				I66x <= 1873;
				I67x <= 1979;
				I68x <= 1896;
				I69x <= 1444;
				I70x <= 1454;
				I71x <= 1088;
				I72x <= 938;
				I73x <= 765;
				I74x <= 971;
				I75x <= 931;
				I76x <= 885;
				I77x <= 801;
				I78x <= 861;
				I79x <= 911;
				I80x <= 888;
				I81x <= 875;
				I82x <= 918;
				I83x <= 1088;
				I84x <= 2568;
				I85x <= 3803;
				I86x <= 6228;
				I87x <= 8192;
				I88x <= 3327;
				I89x <= 712;
				I90x <= 149;
				I91x <= 113;
				I92x <= 622;
				I93x <= 954;
				I94x <= 934;
				I95x <= 1028;
				I96x <= 1078;
				I97x <= 1147;
				I98x <= 1088;
				I99x <= 1194;
				I100x <= 1267;
				I101x <= 1364;
				I102x <= 1354;
				I103x <= 1470;
				I104x <= 1450;
				I105x <= 1620;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111011:begin
				I0x <= 7963;
				I1x <= 7124;
				I2x <= 5138;
				I3x <= 3800;
				I4x <= 1335;
				I5x <= 168;
				I6x <= 518;
				I7x <= 1047;
				I8x <= 2035;
				I9x <= 3314;
				I10x <= 4219;
				I11x <= 4411;
				I12x <= 4504;
				I13x <= 4603;
				I14x <= 4669;
				I15x <= 4685;
				I16x <= 4705;
				I17x <= 4682;
				I18x <= 4692;
				I19x <= 4755;
				I20x <= 4827;
				I21x <= 4781;
				I22x <= 4821;
				I23x <= 4791;
				I24x <= 4844;
				I25x <= 4877;
				I26x <= 4827;
				I27x <= 4788;
				I28x <= 4804;
				I29x <= 4801;
				I30x <= 4785;
				I31x <= 4834;
				I32x <= 4831;
				I33x <= 4794;
				I34x <= 4831;
				I35x <= 4804;
				I36x <= 4808;
				I37x <= 4814;
				I38x <= 4785;
				I39x <= 4712;
				I40x <= 4761;
				I41x <= 4745;
				I42x <= 4745;
				I43x <= 4735;
				I44x <= 4811;
				I45x <= 4821;
				I46x <= 4814;
				I47x <= 4768;
				I48x <= 4765;
				I49x <= 4808;
				I50x <= 4794;
				I51x <= 4768;
				I52x <= 4788;
				I53x <= 4768;
				I54x <= 4781;
				I55x <= 4808;
				I56x <= 4831;
				I57x <= 4864;
				I58x <= 4791;
				I59x <= 4851;
				I60x <= 4785;
				I61x <= 4808;
				I62x <= 4834;
				I63x <= 4775;
				I64x <= 4761;
				I65x <= 4794;
				I66x <= 4738;
				I67x <= 4808;
				I68x <= 4725;
				I69x <= 4808;
				I70x <= 4722;
				I71x <= 4715;
				I72x <= 4708;
				I73x <= 4725;
				I74x <= 4781;
				I75x <= 4742;
				I76x <= 4689;
				I77x <= 4718;
				I78x <= 4692;
				I79x <= 4732;
				I80x <= 4732;
				I81x <= 4732;
				I82x <= 4758;
				I83x <= 4755;
				I84x <= 4689;
				I85x <= 4732;
				I86x <= 4722;
				I87x <= 4695;
				I88x <= 4725;
				I89x <= 4715;
				I90x <= 4765;
				I91x <= 4718;
				I92x <= 4755;
				I93x <= 4682;
				I94x <= 4689;
				I95x <= 4712;
				I96x <= 4705;
				I97x <= 4682;
				I98x <= 4758;
				I99x <= 4728;
				I100x <= 4692;
				I101x <= 4761;
				I102x <= 4758;
				I103x <= 4738;
				I104x <= 4748;
				I105x <= 4732;
				I106x <= 4695;
				I107x <= 4732;
				I108x <= 4689;
				I109x <= 4728;
				I110x <= 4758;
				I111x <= 4801;
				I112x <= 4768;
				I113x <= 4785;
				I114x <= 5019;
				I115x <= 5247;
				I116x <= 5260;
				I117x <= 5277;
				I118x <= 5032;
				I119x <= 5217;
				I120x <= 5082;
				I121x <= 4827;
				I122x <= 4897;
				I123x <= 4976;
				I124x <= 4894;
				I125x <= 4775;
				I126x <= 4599;
				I127x <= 4580;
				I128x <= 4580;
				I129x <= 4530;
				I130x <= 4537;
				I131x <= 4556;
				I132x <= 4563;
				I133x <= 4570;
				I134x <= 4566;
				I135x <= 4560;
				I136x <= 4576;
				I137x <= 4623;
				I138x <= 4632;
				I139x <= 4811;
				I140x <= 5184;
				I141x <= 5492;
				I142x <= 5997;
				I143x <= 7762;
				I144x <= 8192;
				I145x <= 5792;
				I146x <= 3896;
				I147x <= 2052;
				I148x <= 0;
				I149x <= 221;
				I150x <= 713;
				I151x <= 1391;
				I152x <= 2716;
				I153x <= 3978;
				I154x <= 4398;
				I155x <= 4530;
				I156x <= 4599;
				I157x <= 4699;
				I158x <= 4659;
				I159x <= 4738;
				I160x <= 4761;
				I161x <= 4775;
				I162x <= 4801;
				I163x <= 4775;
				I164x <= 4758;
				I165x <= 4748;
				I166x <= 4804;
				I167x <= 4804;
				I168x <= 4761;
				I169x <= 4837;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111100:begin
				I0x <= 8192;
				I1x <= 5333;
				I2x <= 2038;
				I3x <= 233;
				I4x <= 950;
				I5x <= 1459;
				I6x <= 1597;
				I7x <= 1589;
				I8x <= 1688;
				I9x <= 1662;
				I10x <= 1606;
				I11x <= 1589;
				I12x <= 1822;
				I13x <= 1800;
				I14x <= 1882;
				I15x <= 1770;
				I16x <= 1934;
				I17x <= 1826;
				I18x <= 2176;
				I19x <= 1813;
				I20x <= 2029;
				I21x <= 1947;
				I22x <= 2167;
				I23x <= 2154;
				I24x <= 2301;
				I25x <= 2228;
				I26x <= 2435;
				I27x <= 2444;
				I28x <= 2375;
				I29x <= 2474;
				I30x <= 2426;
				I31x <= 2526;
				I32x <= 2508;
				I33x <= 2655;
				I34x <= 2487;
				I35x <= 2202;
				I36x <= 2405;
				I37x <= 2245;
				I38x <= 2392;
				I39x <= 1861;
				I40x <= 1748;
				I41x <= 1943;
				I42x <= 1900;
				I43x <= 1934;
				I44x <= 1917;
				I45x <= 1675;
				I46x <= 1835;
				I47x <= 1835;
				I48x <= 1956;
				I49x <= 1982;
				I50x <= 1774;
				I51x <= 1831;
				I52x <= 1684;
				I53x <= 1731;
				I54x <= 1818;
				I55x <= 1878;
				I56x <= 1973;
				I57x <= 1930;
				I58x <= 1813;
				I59x <= 1891;
				I60x <= 1809;
				I61x <= 1856;
				I62x <= 1666;
				I63x <= 1826;
				I64x <= 1891;
				I65x <= 1567;
				I66x <= 1951;
				I67x <= 1723;
				I68x <= 1705;
				I69x <= 1671;
				I70x <= 1567;
				I71x <= 1822;
				I72x <= 1645;
				I73x <= 1727;
				I74x <= 1800;
				I75x <= 1645;
				I76x <= 1869;
				I77x <= 1515;
				I78x <= 1507;
				I79x <= 1701;
				I80x <= 1740;
				I81x <= 2051;
				I82x <= 2310;
				I83x <= 2245;
				I84x <= 2323;
				I85x <= 2236;
				I86x <= 2254;
				I87x <= 2560;
				I88x <= 2737;
				I89x <= 2413;
				I90x <= 1973;
				I91x <= 1632;
				I92x <= 1351;
				I93x <= 1394;
				I94x <= 1334;
				I95x <= 1377;
				I96x <= 1183;
				I97x <= 1170;
				I98x <= 1075;
				I99x <= 1148;
				I100x <= 1006;
				I101x <= 1049;
				I102x <= 915;
				I103x <= 1429;
				I104x <= 997;
				I105x <= 1312;
				I106x <= 2349;
				I107x <= 4655;
				I108x <= 7643;
				I109x <= 6101;
				I110x <= 2310;
				I111x <= 0;
				I112x <= 462;
				I113x <= 1368;
				I114x <= 1243;
				I115x <= 1334;
				I116x <= 1347;
				I117x <= 1455;
				I118x <= 1485;
				I119x <= 1295;
				I120x <= 1174;
				I121x <= 1399;
				I122x <= 1450;
				I123x <= 1563;
				I124x <= 1351;
				I125x <= 1485;
				I126x <= 1567;
				I127x <= 1472;
				I128x <= 1757;
				I129x <= 1679;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111101:begin
				I0x <= 7848;
				I1x <= 5826;
				I2x <= 581;
				I3x <= 0;
				I4x <= 1044;
				I5x <= 865;
				I6x <= 410;
				I7x <= 529;
				I8x <= 328;
				I9x <= 537;
				I10x <= 395;
				I11x <= 626;
				I12x <= 447;
				I13x <= 276;
				I14x <= 552;
				I15x <= 678;
				I16x <= 701;
				I17x <= 656;
				I18x <= 581;
				I19x <= 872;
				I20x <= 790;
				I21x <= 940;
				I22x <= 1134;
				I23x <= 1208;
				I24x <= 1305;
				I25x <= 1148;
				I26x <= 1328;
				I27x <= 1492;
				I28x <= 1671;
				I29x <= 1984;
				I30x <= 1932;
				I31x <= 1984;
				I32x <= 2059;
				I33x <= 1701;
				I34x <= 1962;
				I35x <= 1738;
				I36x <= 1469;
				I37x <= 1432;
				I38x <= 1216;
				I39x <= 1298;
				I40x <= 1275;
				I41x <= 1290;
				I42x <= 1410;
				I43x <= 1298;
				I44x <= 1305;
				I45x <= 1268;
				I46x <= 1425;
				I47x <= 1171;
				I48x <= 1328;
				I49x <= 1402;
				I50x <= 1126;
				I51x <= 1134;
				I52x <= 1260;
				I53x <= 1365;
				I54x <= 1410;
				I55x <= 1081;
				I56x <= 1305;
				I57x <= 1365;
				I58x <= 1387;
				I59x <= 1328;
				I60x <= 1290;
				I61x <= 1260;
				I62x <= 1328;
				I63x <= 1850;
				I64x <= 2297;
				I65x <= 2536;
				I66x <= 2917;
				I67x <= 3387;
				I68x <= 3126;
				I69x <= 3446;
				I70x <= 3021;
				I71x <= 2536;
				I72x <= 2230;
				I73x <= 1656;
				I74x <= 1290;
				I75x <= 1096;
				I76x <= 1066;
				I77x <= 1044;
				I78x <= 1029;
				I79x <= 1134;
				I80x <= 1007;
				I81x <= 1037;
				I82x <= 813;
				I83x <= 1410;
				I84x <= 3551;
				I85x <= 5476;
				I86x <= 6789;
				I87x <= 8192;
				I88x <= 3797;
				I89x <= 74;
				I90x <= 1738;
				I91x <= 1589;
				I92x <= 1104;
				I93x <= 977;
				I94x <= 1014;
				I95x <= 1044;
				I96x <= 969;
				I97x <= 1074;
				I98x <= 1051;
				I99x <= 1178;
				I100x <= 1044;
				I101x <= 932;
				I102x <= 1044;
				I103x <= 977;
				I104x <= 1134;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111110:begin
				I0x <= 7555;
				I1x <= 5702;
				I2x <= 5104;
				I3x <= 1177;
				I4x <= 1177;
				I5x <= 849;
				I6x <= 0;
				I7x <= 723;
				I8x <= 607;
				I9x <= 501;
				I10x <= 617;
				I11x <= 723;
				I12x <= 771;
				I13x <= 578;
				I14x <= 810;
				I15x <= 926;
				I16x <= 897;
				I17x <= 742;
				I18x <= 1022;
				I19x <= 1167;
				I20x <= 1080;
				I21x <= 1331;
				I22x <= 1717;
				I23x <= 1437;
				I24x <= 1958;
				I25x <= 2161;
				I26x <= 2113;
				I27x <= 2566;
				I28x <= 2267;
				I29x <= 2151;
				I30x <= 1823;
				I31x <= 1978;
				I32x <= 1939;
				I33x <= 1678;
				I34x <= 1842;
				I35x <= 1630;
				I36x <= 1264;
				I37x <= 1350;
				I38x <= 1447;
				I39x <= 1235;
				I40x <= 955;
				I41x <= 1090;
				I42x <= 1264;
				I43x <= 1022;
				I44x <= 1514;
				I45x <= 1312;
				I46x <= 1399;
				I47x <= 1341;
				I48x <= 1495;
				I49x <= 1678;
				I50x <= 1399;
				I51x <= 1302;
				I52x <= 1871;
				I53x <= 1321;
				I54x <= 1466;
				I55x <= 1756;
				I56x <= 1466;
				I57x <= 1495;
				I58x <= 1292;
				I59x <= 1553;
				I60x <= 1321;
				I61x <= 1302;
				I62x <= 1592;
				I63x <= 1553;
				I64x <= 1437;
				I65x <= 2026;
				I66x <= 1823;
				I67x <= 1717;
				I68x <= 1640;
				I69x <= 1495;
				I70x <= 1958;
				I71x <= 1968;
				I72x <= 2711;
				I73x <= 2981;
				I74x <= 2749;
				I75x <= 3406;
				I76x <= 4120;
				I77x <= 4457;
				I78x <= 3579;
				I79x <= 2875;
				I80x <= 2450;
				I81x <= 2499;
				I82x <= 2470;
				I83x <= 2084;
				I84x <= 1910;
				I85x <= 1785;
				I86x <= 2171;
				I87x <= 2605;
				I88x <= 2402;
				I89x <= 2122;
				I90x <= 3801;
				I91x <= 6320;
				I92x <= 7632;
				I93x <= 8192;
				I94x <= 6358;
				I95x <= 4920;
				I96x <= 1939;
				I97x <= 2209;
				I98x <= 2084;
				I99x <= 1736;
				I100x <= 1505;
				I101x <= 1862;
				I102x <= 1746;
				I103x <= 1659;
				I104x <= 2257;
				I105x <= 1939;
				I106x <= 2209;
				I107x <= 2180;
				I108x <= 2364;
				I109x <= 2392;
				I110x <= 2161;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b00111111:begin
				I0x <= 8192;
				I1x <= 6032;
				I2x <= 3767;
				I3x <= 3141;
				I4x <= 2224;
				I5x <= 966;
				I6x <= 657;
				I7x <= 374;
				I8x <= 460;
				I9x <= 230;
				I10x <= 444;
				I11x <= 374;
				I12x <= 345;
				I13x <= 477;
				I14x <= 287;
				I15x <= 472;
				I16x <= 444;
				I17x <= 493;
				I18x <= 575;
				I19x <= 366;
				I20x <= 641;
				I21x <= 620;
				I22x <= 699;
				I23x <= 773;
				I24x <= 649;
				I25x <= 904;
				I26x <= 937;
				I27x <= 1032;
				I28x <= 1225;
				I29x <= 1200;
				I30x <= 1603;
				I31x <= 1801;
				I32x <= 2068;
				I33x <= 2422;
				I34x <= 2434;
				I35x <= 2808;
				I36x <= 2952;
				I37x <= 3067;
				I38x <= 3059;
				I39x <= 2644;
				I40x <= 2529;
				I41x <= 2224;
				I42x <= 1957;
				I43x <= 1747;
				I44x <= 1332;
				I45x <= 1328;
				I46x <= 1217;
				I47x <= 1135;
				I48x <= 1126;
				I49x <= 908;
				I50x <= 1126;
				I51x <= 1081;
				I52x <= 1089;
				I53x <= 1102;
				I54x <= 888;
				I55x <= 1110;
				I56x <= 1048;
				I57x <= 1089;
				I58x <= 1114;
				I59x <= 945;
				I60x <= 1093;
				I61x <= 1028;
				I62x <= 1052;
				I63x <= 1093;
				I64x <= 875;
				I65x <= 1089;
				I66x <= 1044;
				I67x <= 1019;
				I68x <= 1015;
				I69x <= 810;
				I70x <= 1032;
				I71x <= 954;
				I72x <= 991;
				I73x <= 904;
				I74x <= 773;
				I75x <= 970;
				I76x <= 949;
				I77x <= 982;
				I78x <= 871;
				I79x <= 760;
				I80x <= 1007;
				I81x <= 945;
				I82x <= 921;
				I83x <= 896;
				I84x <= 773;
				I85x <= 1122;
				I86x <= 1213;
				I87x <= 1250;
				I88x <= 1402;
				I89x <= 1221;
				I90x <= 1402;
				I91x <= 1468;
				I92x <= 1472;
				I93x <= 1287;
				I94x <= 1246;
				I95x <= 1299;
				I96x <= 1114;
				I97x <= 991;
				I98x <= 1003;
				I99x <= 674;
				I100x <= 760;
				I101x <= 620;
				I102x <= 653;
				I103x <= 583;
				I104x <= 756;
				I105x <= 1677;
				I106x <= 2817;
				I107x <= 5136;
				I108x <= 8093;
				I109x <= 5436;
				I110x <= 3326;
				I111x <= 2467;
				I112x <= 1517;
				I113x <= 699;
				I114x <= 333;
				I115x <= 407;
				I116x <= 168;
				I117x <= 189;
				I118x <= 205;
				I119x <= 98;
				I120x <= 267;
				I121x <= 176;
				I122x <= 135;
				I123x <= 180;
				I124x <= 0;
				I125x <= 238;
				I126x <= 238;
				I127x <= 213;
				I128x <= 259;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000000:begin
				I0x <= 8192;
				I1x <= 6119;
				I2x <= 3068;
				I3x <= 1628;
				I4x <= 1952;
				I5x <= 1460;
				I6x <= 715;
				I7x <= 573;
				I8x <= 586;
				I9x <= 547;
				I10x <= 400;
				I11x <= 892;
				I12x <= 633;
				I13x <= 801;
				I14x <= 857;
				I15x <= 736;
				I16x <= 900;
				I17x <= 810;
				I18x <= 719;
				I19x <= 590;
				I20x <= 672;
				I21x <= 736;
				I22x <= 555;
				I23x <= 551;
				I24x <= 564;
				I25x <= 581;
				I26x <= 655;
				I27x <= 965;
				I28x <= 836;
				I29x <= 848;
				I30x <= 818;
				I31x <= 1271;
				I32x <= 1159;
				I33x <= 1141;
				I34x <= 1103;
				I35x <= 1133;
				I36x <= 1249;
				I37x <= 1146;
				I38x <= 1245;
				I39x <= 1258;
				I40x <= 1297;
				I41x <= 1417;
				I42x <= 1327;
				I43x <= 1529;
				I44x <= 1391;
				I45x <= 1210;
				I46x <= 1422;
				I47x <= 1594;
				I48x <= 1607;
				I49x <= 1861;
				I50x <= 1891;
				I51x <= 1887;
				I52x <= 1637;
				I53x <= 1581;
				I54x <= 1615;
				I55x <= 1366;
				I56x <= 1482;
				I57x <= 1396;
				I58x <= 1163;
				I59x <= 913;
				I60x <= 848;
				I61x <= 792;
				I62x <= 1034;
				I63x <= 801;
				I64x <= 853;
				I65x <= 0;
				I66x <= 517;
				I67x <= 495;
				I68x <= 418;
				I69x <= 2745;
				I70x <= 7502;
				I71x <= 7765;
				I72x <= 5434;
				I73x <= 2658;
				I74x <= 1771;
				I75x <= 1689;
				I76x <= 1146;
				I77x <= 693;
				I78x <= 741;
				I79x <= 560;
				I80x <= 594;
				I81x <= 564;
				I82x <= 693;
				I83x <= 633;
				I84x <= 719;
				I85x <= 0;
				I86x <= 0;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000001:begin
				I0x <= 8164;
				I1x <= 6251;
				I2x <= 2041;
				I3x <= 827;
				I4x <= 372;
				I5x <= 952;
				I6x <= 1328;
				I7x <= 1418;
				I8x <= 1609;
				I9x <= 1585;
				I10x <= 1589;
				I11x <= 1655;
				I12x <= 1703;
				I13x <= 1832;
				I14x <= 1870;
				I15x <= 1724;
				I16x <= 1915;
				I17x <= 1940;
				I18x <= 2141;
				I19x <= 2127;
				I20x <= 2183;
				I21x <= 2322;
				I22x <= 2430;
				I23x <= 2256;
				I24x <= 2510;
				I25x <= 2496;
				I26x <= 2670;
				I27x <= 2680;
				I28x <= 2771;
				I29x <= 2746;
				I30x <= 2527;
				I31x <= 2430;
				I32x <= 2315;
				I33x <= 2253;
				I34x <= 2228;
				I35x <= 1908;
				I36x <= 1884;
				I37x <= 1571;
				I38x <= 1769;
				I39x <= 1686;
				I40x <= 1592;
				I41x <= 1748;
				I42x <= 1554;
				I43x <= 1648;
				I44x <= 1543;
				I45x <= 1787;
				I46x <= 1717;
				I47x <= 1863;
				I48x <= 1867;
				I49x <= 1846;
				I50x <= 1908;
				I51x <= 1961;
				I52x <= 1745;
				I53x <= 1815;
				I54x <= 1679;
				I55x <= 1665;
				I56x <= 1696;
				I57x <= 1522;
				I58x <= 1682;
				I59x <= 1540;
				I60x <= 1505;
				I61x <= 1627;
				I62x <= 1509;
				I63x <= 1644;
				I64x <= 1665;
				I65x <= 1849;
				I66x <= 2114;
				I67x <= 2065;
				I68x <= 1981;
				I69x <= 2211;
				I70x <= 2162;
				I71x <= 2127;
				I72x <= 1710;
				I73x <= 1735;
				I74x <= 1540;
				I75x <= 1185;
				I76x <= 1227;
				I77x <= 1168;
				I78x <= 1210;
				I79x <= 1189;
				I80x <= 1164;
				I81x <= 1164;
				I82x <= 1112;
				I83x <= 1230;
				I84x <= 1237;
				I85x <= 1105;
				I86x <= 1192;
				I87x <= 2632;
				I88x <= 3657;
				I89x <= 6276;
				I90x <= 8192;
				I91x <= 4829;
				I92x <= 945;
				I93x <= 344;
				I94x <= 0;
				I95x <= 531;
				I96x <= 931;
				I97x <= 1112;
				I98x <= 1060;
				I99x <= 1251;
				I100x <= 1199;
				I101x <= 1296;
				I102x <= 1241;
				I103x <= 1460;
				I104x <= 1474;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000010:begin
				I0x <= 7452;
				I1x <= 3027;
				I2x <= 0;
				I3x <= 121;
				I4x <= 1154;
				I5x <= 1225;
				I6x <= 1113;
				I7x <= 718;
				I8x <= 1144;
				I9x <= 1174;
				I10x <= 1022;
				I11x <= 1154;
				I12x <= 1539;
				I13x <= 840;
				I14x <= 1579;
				I15x <= 1741;
				I16x <= 1194;
				I17x <= 1458;
				I18x <= 1630;
				I19x <= 1842;
				I20x <= 2045;
				I21x <= 1751;
				I22x <= 2106;
				I23x <= 2379;
				I24x <= 2572;
				I25x <= 2420;
				I26x <= 2268;
				I27x <= 2653;
				I28x <= 1964;
				I29x <= 1812;
				I30x <= 2085;
				I31x <= 1883;
				I32x <= 1913;
				I33x <= 1458;
				I34x <= 1954;
				I35x <= 1205;
				I36x <= 1377;
				I37x <= 1397;
				I38x <= 1377;
				I39x <= 1539;
				I40x <= 1397;
				I41x <= 1488;
				I42x <= 1518;
				I43x <= 1488;
				I44x <= 1934;
				I45x <= 1842;
				I46x <= 1448;
				I47x <= 1680;
				I48x <= 1853;
				I49x <= 2015;
				I50x <= 1772;
				I51x <= 1761;
				I52x <= 1923;
				I53x <= 1934;
				I54x <= 1660;
				I55x <= 1873;
				I56x <= 1741;
				I57x <= 1367;
				I58x <= 2065;
				I59x <= 1731;
				I60x <= 1468;
				I61x <= 1417;
				I62x <= 1761;
				I63x <= 2328;
				I64x <= 2592;
				I65x <= 2956;
				I66x <= 3706;
				I67x <= 2369;
				I68x <= 3584;
				I69x <= 3250;
				I70x <= 2470;
				I71x <= 2713;
				I72x <= 2339;
				I73x <= 1670;
				I74x <= 1215;
				I75x <= 1073;
				I76x <= 820;
				I77x <= 911;
				I78x <= 1093;
				I79x <= 577;
				I80x <= 951;
				I81x <= 384;
				I82x <= 860;
				I83x <= 2258;
				I84x <= 2622;
				I85x <= 2946;
				I86x <= 5781;
				I87x <= 8192;
				I88x <= 5387;
				I89x <= 1397;
				I90x <= 313;
				I91x <= 1437;
				I92x <= 1316;
				I93x <= 840;
				I94x <= 1468;
				I95x <= 1367;
				I96x <= 1316;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000011:begin
				I0x <= 7928;
				I1x <= 5483;
				I2x <= 2147;
				I3x <= 1083;
				I4x <= 116;
				I5x <= 37;
				I6x <= 101;
				I7x <= 41;
				I8x <= 33;
				I9x <= 26;
				I10x <= 82;
				I11x <= 116;
				I12x <= 157;
				I13x <= 176;
				I14x <= 112;
				I15x <= 161;
				I16x <= 195;
				I17x <= 188;
				I18x <= 240;
				I19x <= 173;
				I20x <= 195;
				I21x <= 161;
				I22x <= 127;
				I23x <= 124;
				I24x <= 0;
				I25x <= 229;
				I26x <= 240;
				I27x <= 173;
				I28x <= 289;
				I29x <= 297;
				I30x <= 440;
				I31x <= 511;
				I32x <= 552;
				I33x <= 699;
				I34x <= 748;
				I35x <= 1000;
				I36x <= 1120;
				I37x <= 1143;
				I38x <= 1286;
				I39x <= 1256;
				I40x <= 1241;
				I41x <= 1143;
				I42x <= 992;
				I43x <= 940;
				I44x <= 906;
				I45x <= 940;
				I46x <= 929;
				I47x <= 940;
				I48x <= 944;
				I49x <= 846;
				I50x <= 842;
				I51x <= 865;
				I52x <= 789;
				I53x <= 940;
				I54x <= 819;
				I55x <= 883;
				I56x <= 974;
				I57x <= 981;
				I58x <= 1154;
				I59x <= 1113;
				I60x <= 1132;
				I61x <= 1147;
				I62x <= 1071;
				I63x <= 1165;
				I64x <= 1143;
				I65x <= 1177;
				I66x <= 1109;
				I67x <= 1150;
				I68x <= 1184;
				I69x <= 1053;
				I70x <= 1147;
				I71x <= 1147;
				I72x <= 1102;
				I73x <= 1271;
				I74x <= 1241;
				I75x <= 1391;
				I76x <= 1308;
				I77x <= 1305;
				I78x <= 1489;
				I79x <= 1402;
				I80x <= 1527;
				I81x <= 1448;
				I82x <= 1433;
				I83x <= 1515;
				I84x <= 1455;
				I85x <= 1448;
				I86x <= 1399;
				I87x <= 1440;
				I88x <= 1463;
				I89x <= 1361;
				I90x <= 1448;
				I91x <= 1575;
				I92x <= 1718;
				I93x <= 2027;
				I94x <= 1903;
				I95x <= 1982;
				I96x <= 2132;
				I97x <= 2061;
				I98x <= 2128;
				I99x <= 2110;
				I100x <= 1786;
				I101x <= 1538;
				I102x <= 1214;
				I103x <= 1079;
				I104x <= 1090;
				I105x <= 1038;
				I106x <= 1109;
				I107x <= 1045;
				I108x <= 1120;
				I109x <= 816;
				I110x <= 154;
				I111x <= 214;
				I112x <= 2561;
				I113x <= 6574;
				I114x <= 8192;
				I115x <= 6021;
				I116x <= 3302;
				I117x <= 2313;
				I118x <= 1339;
				I119x <= 921;
				I120x <= 917;
				I121x <= 944;
				I122x <= 834;
				I123x <= 876;
				I124x <= 857;
				I125x <= 827;
				I126x <= 910;
				I127x <= 744;
				I128x <= 898;
				I129x <= 804;
				I130x <= 940;
				I131x <= 865;
				I132x <= 767;
				I133x <= 913;
				I134x <= 898;
				I135x <= 977;
				I136x <= 940;
				I137x <= 977;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000100:begin
				I0x <= 8192;
				I1x <= 3607;
				I2x <= 2546;
				I3x <= 307;
				I4x <= 44;
				I5x <= 0;
				I6x <= 1960;
				I7x <= 2323;
				I8x <= 2378;
				I9x <= 2747;
				I10x <= 2596;
				I11x <= 2758;
				I12x <= 3048;
				I13x <= 2780;
				I14x <= 2903;
				I15x <= 3043;
				I16x <= 2981;
				I17x <= 3115;
				I18x <= 2987;
				I19x <= 3127;
				I20x <= 3216;
				I21x <= 3277;
				I22x <= 3395;
				I23x <= 3322;
				I24x <= 3255;
				I25x <= 3149;
				I26x <= 3311;
				I27x <= 3473;
				I28x <= 3585;
				I29x <= 3735;
				I30x <= 3501;
				I31x <= 3568;
				I32x <= 4054;
				I33x <= 3797;
				I34x <= 3791;
				I35x <= 3808;
				I36x <= 3864;
				I37x <= 3579;
				I38x <= 3445;
				I39x <= 3166;
				I40x <= 2685;
				I41x <= 2769;
				I42x <= 2646;
				I43x <= 2753;
				I44x <= 2747;
				I45x <= 2702;
				I46x <= 2658;
				I47x <= 2658;
				I48x <= 3009;
				I49x <= 2820;
				I50x <= 2792;
				I51x <= 3182;
				I52x <= 3160;
				I53x <= 3060;
				I54x <= 3512;
				I55x <= 3233;
				I56x <= 3171;
				I57x <= 3261;
				I58x <= 3194;
				I59x <= 2948;
				I60x <= 3333;
				I61x <= 3004;
				I62x <= 2808;
				I63x <= 3255;
				I64x <= 3182;
				I65x <= 2903;
				I66x <= 3015;
				I67x <= 3043;
				I68x <= 3143;
				I69x <= 3088;
				I70x <= 3021;
				I71x <= 3099;
				I72x <= 3093;
				I73x <= 2998;
				I74x <= 2948;
				I75x <= 3182;
				I76x <= 2898;
				I77x <= 2998;
				I78x <= 2920;
				I79x <= 3300;
				I80x <= 2993;
				I81x <= 2954;
				I82x <= 2613;
				I83x <= 2903;
				I84x <= 3266;
				I85x <= 3255;
				I86x <= 3093;
				I87x <= 2998;
				I88x <= 3082;
				I89x <= 3210;
				I90x <= 3060;
				I91x <= 2847;
				I92x <= 3071;
				I93x <= 2909;
				I94x <= 3021;
				I95x <= 3177;
				I96x <= 3261;
				I97x <= 3071;
				I98x <= 3048;
				I99x <= 3132;
				I100x <= 3266;
				I101x <= 3618;
				I102x <= 3378;
				I103x <= 3601;
				I104x <= 3998;
				I105x <= 4551;
				I106x <= 4422;
				I107x <= 4327;
				I108x <= 3981;
				I109x <= 3707;
				I110x <= 3367;
				I111x <= 3071;
				I112x <= 2898;
				I113x <= 2842;
				I114x <= 3060;
				I115x <= 2920;
				I116x <= 2909;
				I117x <= 3015;
				I118x <= 3847;
				I119x <= 4590;
				I120x <= 6282;
				I121x <= 7990;
				I122x <= 6756;
				I123x <= 3166;
				I124x <= 1569;
				I125x <= 301;
				I126x <= 374;
				I127x <= 1429;
				I128x <= 2959;
				I129x <= 2875;
				I130x <= 3333;
				I131x <= 2970;
				I132x <= 3652;
				I133x <= 3384;
				I134x <= 3478;
				I135x <= 3540;
				I136x <= 3400;
				I137x <= 3741;
				I138x <= 3266;
				I139x <= 3668;
				I140x <= 3646;
				I141x <= 3523;
				I142x <= 3903;
				I143x <= 3551;
				I144x <= 3702;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000101:begin
				I0x <= 7982;
				I1x <= 4537;
				I2x <= 16;
				I3x <= 511;
				I4x <= 1603;
				I5x <= 1087;
				I6x <= 1194;
				I7x <= 995;
				I8x <= 1124;
				I9x <= 1248;
				I10x <= 1221;
				I11x <= 1394;
				I12x <= 979;
				I13x <= 1340;
				I14x <= 1302;
				I15x <= 1275;
				I16x <= 1577;
				I17x <= 1286;
				I18x <= 1420;
				I19x <= 1523;
				I20x <= 1453;
				I21x <= 1587;
				I22x <= 1281;
				I23x <= 1340;
				I24x <= 1324;
				I25x <= 1178;
				I26x <= 1603;
				I27x <= 1286;
				I28x <= 1410;
				I29x <= 1431;
				I30x <= 1754;
				I31x <= 1743;
				I32x <= 1593;
				I33x <= 1733;
				I34x <= 1657;
				I35x <= 1813;
				I36x <= 1959;
				I37x <= 1603;
				I38x <= 1910;
				I39x <= 1840;
				I40x <= 1851;
				I41x <= 1937;
				I42x <= 1523;
				I43x <= 1652;
				I44x <= 1603;
				I45x <= 1630;
				I46x <= 1706;
				I47x <= 1566;
				I48x <= 1851;
				I49x <= 1711;
				I50x <= 1878;
				I51x <= 1964;
				I52x <= 1614;
				I53x <= 1943;
				I54x <= 2115;
				I55x <= 2572;
				I56x <= 3024;
				I57x <= 2610;
				I58x <= 2884;
				I59x <= 2814;
				I60x <= 3396;
				I61x <= 3487;
				I62x <= 2260;
				I63x <= 2196;
				I64x <= 1846;
				I65x <= 1603;
				I66x <= 1711;
				I67x <= 1297;
				I68x <= 1496;
				I69x <= 1496;
				I70x <= 1464;
				I71x <= 1743;
				I72x <= 1345;
				I73x <= 974;
				I74x <= 710;
				I75x <= 2761;
				I76x <= 5366;
				I77x <= 8192;
				I78x <= 5533;
				I79x <= 1146;
				I80x <= 0;
				I81x <= 1695;
				I82x <= 1114;
				I83x <= 1340;
				I84x <= 1189;
				I85x <= 1189;
				I86x <= 1377;
				I87x <= 979;
				I88x <= 1286;
				I89x <= 1167;
				I90x <= 1194;
				I91x <= 1350;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000110:begin
				I0x <= 8192;
				I1x <= 2447;
				I2x <= 725;
				I3x <= 184;
				I4x <= 620;
				I5x <= 2150;
				I6x <= 2315;
				I7x <= 2051;
				I8x <= 2473;
				I9x <= 1998;
				I10x <= 2552;
				I11x <= 2394;
				I12x <= 2420;
				I13x <= 2882;
				I14x <= 2440;
				I15x <= 2829;
				I16x <= 2823;
				I17x <= 2611;
				I18x <= 3350;
				I19x <= 3007;
				I20x <= 3436;
				I21x <= 3634;
				I22x <= 3772;
				I23x <= 4504;
				I24x <= 4379;
				I25x <= 5006;
				I26x <= 5223;
				I27x <= 5421;
				I28x <= 6028;
				I29x <= 5672;
				I30x <= 5923;
				I31x <= 5731;
				I32x <= 5032;
				I33x <= 5032;
				I34x <= 4016;
				I35x <= 3818;
				I36x <= 3324;
				I37x <= 2823;
				I38x <= 2908;
				I39x <= 2361;
				I40x <= 2658;
				I41x <= 2460;
				I42x <= 2176;
				I43x <= 2552;
				I44x <= 2031;
				I45x <= 2552;
				I46x <= 2295;
				I47x <= 2104;
				I48x <= 2605;
				I49x <= 2071;
				I50x <= 2466;
				I51x <= 2315;
				I52x <= 2084;
				I53x <= 2394;
				I54x <= 1919;
				I55x <= 2196;
				I56x <= 2137;
				I57x <= 1892;
				I58x <= 2295;
				I59x <= 1701;
				I60x <= 1998;
				I61x <= 1925;
				I62x <= 1794;
				I63x <= 2064;
				I64x <= 1681;
				I65x <= 1932;
				I66x <= 1807;
				I67x <= 2235;
				I68x <= 3106;
				I69x <= 2730;
				I70x <= 2994;
				I71x <= 3139;
				I72x <= 2770;
				I73x <= 2809;
				I74x <= 2044;
				I75x <= 2354;
				I76x <= 2123;
				I77x <= 1701;
				I78x <= 1932;
				I79x <= 1418;
				I80x <= 1721;
				I81x <= 1444;
				I82x <= 1470;
				I83x <= 1807;
				I84x <= 1160;
				I85x <= 1767;
				I86x <= 2783;
				I87x <= 1741;
				I88x <= 8013;
				I89x <= 5461;
				I90x <= 1240;
				I91x <= 310;
				I92x <= 0;
				I93x <= 1668;
				I94x <= 1662;
				I95x <= 1985;
				I96x <= 1925;
				I97x <= 1714;
				I98x <= 2143;
				I99x <= 1728;
				I100x <= 2130;
				I101x <= 2117;
				I102x <= 2110;
				I103x <= 2625;
				I104x <= 2143;
				I105x <= 2565;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01000111:begin
				I0x <= 8192;
				I1x <= 6837;
				I2x <= 6284;
				I3x <= 5376;
				I4x <= 4261;
				I5x <= 3768;
				I6x <= 3217;
				I7x <= 2425;
				I8x <= 2083;
				I9x <= 2392;
				I10x <= 2601;
				I11x <= 1921;
				I12x <= 2675;
				I13x <= 2160;
				I14x <= 2441;
				I15x <= 2309;
				I16x <= 2224;
				I17x <= 2270;
				I18x <= 2138;
				I19x <= 2956;
				I20x <= 2573;
				I21x <= 2281;
				I22x <= 2565;
				I23x <= 2535;
				I24x <= 2573;
				I25x <= 2210;
				I26x <= 2639;
				I27x <= 2529;
				I28x <= 3116;
				I29x <= 2392;
				I30x <= 2678;
				I31x <= 2697;
				I32x <= 2359;
				I33x <= 2521;
				I34x <= 2645;
				I35x <= 2441;
				I36x <= 2937;
				I37x <= 2997;
				I38x <= 2901;
				I39x <= 2554;
				I40x <= 2416;
				I41x <= 2893;
				I42x <= 2661;
				I43x <= 2339;
				I44x <= 2807;
				I45x <= 2507;
				I46x <= 2364;
				I47x <= 2507;
				I48x <= 2956;
				I49x <= 2584;
				I50x <= 2458;
				I51x <= 2438;
				I52x <= 2381;
				I53x <= 2521;
				I54x <= 2235;
				I55x <= 2807;
				I56x <= 2491;
				I57x <= 2634;
				I58x <= 2725;
				I59x <= 3157;
				I60x <= 2854;
				I61x <= 3300;
				I62x <= 3446;
				I63x <= 3740;
				I64x <= 3595;
				I65x <= 3556;
				I66x <= 3416;
				I67x <= 3124;
				I68x <= 2857;
				I69x <= 2719;
				I70x <= 2471;
				I71x <= 2392;
				I72x <= 2204;
				I73x <= 2312;
				I74x <= 2078;
				I75x <= 2034;
				I76x <= 1957;
				I77x <= 806;
				I78x <= 0;
				I79x <= 756;
				I80x <= 4398;
				I81x <= 7459;
				I82x <= 8169;
				I83x <= 6947;
				I84x <= 5645;
				I85x <= 5108;
				I86x <= 4291;
				I87x <= 3705;
				I88x <= 2994;
				I89x <= 2281;
				I90x <= 2210;
				I91x <= 2411;
				I92x <= 2254;
				I93x <= 2138;
				I94x <= 2158;
				I95x <= 2166;
				I96x <= 1957;
				I97x <= 2191;
				I98x <= 2111;
				I99x <= 2804;
				I100x <= 2295;
				I101x <= 2048;
				I102x <= 2202;
				I103x <= 2207;
				I104x <= 2226;
				I105x <= 2262;
				I106x <= 2130;
				I107x <= 2083;
				I108x <= 2281;
				I109x <= 2221;
				I110x <= 2224;
				I111x <= 2295;
				I112x <= 2199;
				I113x <= 2028;
				I114x <= 2507;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001000:begin
				I0x <= 7648;
				I1x <= 6438;
				I2x <= 5820;
				I3x <= 5199;
				I4x <= 4254;
				I5x <= 3713;
				I6x <= 3302;
				I7x <= 2653;
				I8x <= 2219;
				I9x <= 2581;
				I10x <= 2129;
				I11x <= 2230;
				I12x <= 2075;
				I13x <= 2101;
				I14x <= 2098;
				I15x <= 2167;
				I16x <= 2244;
				I17x <= 2155;
				I18x <= 2230;
				I19x <= 2086;
				I20x <= 2400;
				I21x <= 2069;
				I22x <= 2083;
				I23x <= 2256;
				I24x <= 2299;
				I25x <= 2276;
				I26x <= 2250;
				I27x <= 2420;
				I28x <= 2316;
				I29x <= 2385;
				I30x <= 2345;
				I31x <= 2259;
				I32x <= 2397;
				I33x <= 2492;
				I34x <= 2351;
				I35x <= 2362;
				I36x <= 2351;
				I37x <= 2362;
				I38x <= 2532;
				I39x <= 2489;
				I40x <= 2348;
				I41x <= 2144;
				I42x <= 2397;
				I43x <= 2316;
				I44x <= 2440;
				I45x <= 2247;
				I46x <= 2336;
				I47x <= 2244;
				I48x <= 2132;
				I49x <= 2187;
				I50x <= 2250;
				I51x <= 1957;
				I52x <= 2356;
				I53x <= 2434;
				I54x <= 2196;
				I55x <= 2299;
				I56x <= 2480;
				I57x <= 2230;
				I58x <= 1761;
				I59x <= 2722;
				I60x <= 2267;
				I61x <= 2147;
				I62x <= 2296;
				I63x <= 2164;
				I64x <= 2345;
				I65x <= 2759;
				I66x <= 2630;
				I67x <= 2753;
				I68x <= 2687;
				I69x <= 2920;
				I70x <= 3138;
				I71x <= 2992;
				I72x <= 3250;
				I73x <= 3299;
				I74x <= 2693;
				I75x <= 2348;
				I76x <= 2020;
				I77x <= 2072;
				I78x <= 1885;
				I79x <= 1902;
				I80x <= 1675;
				I81x <= 1980;
				I82x <= 1991;
				I83x <= 1649;
				I84x <= 640;
				I85x <= 0;
				I86x <= 799;
				I87x <= 3489;
				I88x <= 6789;
				I89x <= 8192;
				I90x <= 6496;
				I91x <= 5352;
				I92x <= 5001;
				I93x <= 3952;
				I94x <= 3584;
				I95x <= 2842;
				I96x <= 1888;
				I97x <= 2299;
				I98x <= 1629;
				I99x <= 1928;
				I100x <= 2104;
				I101x <= 1908;
				I102x <= 1911;
				I103x <= 1876;
				I104x <= 1911;
				I105x <= 1871;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001001:begin
				I0x <= 8192;
				I1x <= 8034;
				I2x <= 4899;
				I3x <= 3435;
				I4x <= 2485;
				I5x <= 2018;
				I6x <= 2313;
				I7x <= 2228;
				I8x <= 2213;
				I9x <= 2142;
				I10x <= 2213;
				I11x <= 2352;
				I12x <= 2328;
				I13x <= 2418;
				I14x <= 2380;
				I15x <= 2399;
				I16x <= 2485;
				I17x <= 2509;
				I18x <= 2595;
				I19x <= 2585;
				I20x <= 2538;
				I21x <= 2709;
				I22x <= 2581;
				I23x <= 2581;
				I24x <= 2523;
				I25x <= 2504;
				I26x <= 2232;
				I27x <= 2299;
				I28x <= 2347;
				I29x <= 2266;
				I30x <= 2180;
				I31x <= 2209;
				I32x <= 2132;
				I33x <= 2170;
				I34x <= 2218;
				I35x <= 2337;
				I36x <= 2576;
				I37x <= 2605;
				I38x <= 2705;
				I39x <= 2638;
				I40x <= 2695;
				I41x <= 2824;
				I42x <= 2748;
				I43x <= 2872;
				I44x <= 2729;
				I45x <= 2814;
				I46x <= 2891;
				I47x <= 2805;
				I48x <= 2848;
				I49x <= 2748;
				I50x <= 2767;
				I51x <= 2781;
				I52x <= 2652;
				I53x <= 2800;
				I54x <= 2676;
				I55x <= 2695;
				I56x <= 2724;
				I57x <= 2614;
				I58x <= 2686;
				I59x <= 2624;
				I60x <= 2667;
				I61x <= 2638;
				I62x <= 2514;
				I63x <= 2614;
				I64x <= 2752;
				I65x <= 3015;
				I66x <= 3292;
				I67x <= 3420;
				I68x <= 3840;
				I69x <= 3979;
				I70x <= 3616;
				I71x <= 3330;
				I72x <= 3067;
				I73x <= 2786;
				I74x <= 2480;
				I75x <= 2356;
				I76x <= 2347;
				I77x <= 2213;
				I78x <= 2342;
				I79x <= 2247;
				I80x <= 1688;
				I81x <= 415;
				I82x <= 0;
				I83x <= 3210;
				I84x <= 6784;
				I85x <= 7948;
				I86x <= 6832;
				I87x <= 3587;
				I88x <= 3048;
				I89x <= 2228;
				I90x <= 2304;
				I91x <= 2275;
				I92x <= 2166;
				I93x <= 2199;
				I94x <= 2175;
				I95x <= 2218;
				I96x <= 2337;
				I97x <= 2323;
				I98x <= 2504;
				I99x <= 2423;
				I100x <= 2495;
				I101x <= 2504;
				I102x <= 2361;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001010:begin
				I0x <= 7886;
				I1x <= 2464;
				I2x <= 686;
				I3x <= 653;
				I4x <= 797;
				I5x <= 867;
				I6x <= 869;
				I7x <= 852;
				I8x <= 810;
				I9x <= 782;
				I10x <= 889;
				I11x <= 767;
				I12x <= 745;
				I13x <= 681;
				I14x <= 701;
				I15x <= 688;
				I16x <= 636;
				I17x <= 722;
				I18x <= 690;
				I19x <= 653;
				I20x <= 743;
				I21x <= 775;
				I22x <= 837;
				I23x <= 914;
				I24x <= 998;
				I25x <= 1162;
				I26x <= 1188;
				I27x <= 1340;
				I28x <= 1372;
				I29x <= 1416;
				I30x <= 1528;
				I31x <= 1472;
				I32x <= 1536;
				I33x <= 1581;
				I34x <= 1534;
				I35x <= 1613;
				I36x <= 1566;
				I37x <= 1515;
				I38x <= 1530;
				I39x <= 1515;
				I40x <= 1568;
				I41x <= 1517;
				I42x <= 1540;
				I43x <= 1555;
				I44x <= 1487;
				I45x <= 1500;
				I46x <= 1416;
				I47x <= 1459;
				I48x <= 1421;
				I49x <= 1404;
				I50x <= 1446;
				I51x <= 1389;
				I52x <= 1421;
				I53x <= 1431;
				I54x <= 1395;
				I55x <= 1451;
				I56x <= 1404;
				I57x <= 1429;
				I58x <= 1446;
				I59x <= 1455;
				I60x <= 1763;
				I61x <= 1846;
				I62x <= 1961;
				I63x <= 1947;
				I64x <= 1797;
				I65x <= 1889;
				I66x <= 1782;
				I67x <= 1711;
				I68x <= 1496;
				I69x <= 1372;
				I70x <= 1380;
				I71x <= 1506;
				I72x <= 1402;
				I73x <= 1348;
				I74x <= 1318;
				I75x <= 1372;
				I76x <= 1316;
				I77x <= 1369;
				I78x <= 1425;
				I79x <= 1361;
				I80x <= 1077;
				I81x <= 592;
				I82x <= 0;
				I83x <= 583;
				I84x <= 3812;
				I85x <= 8192;
				I86x <= 5358;
				I87x <= 1081;
				I88x <= 600;
				I89x <= 718;
				I90x <= 886;
				I91x <= 869;
				I92x <= 850;
				I93x <= 857;
				I94x <= 799;
				I95x <= 854;
				I96x <= 786;
				I97x <= 767;
				I98x <= 760;
				I99x <= 722;
				I100x <= 788;
				I101x <= 701;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001011:begin
				I0x <= 8192;
				I1x <= 8086;
				I2x <= 1422;
				I3x <= 0;
				I4x <= 1151;
				I5x <= 857;
				I6x <= 1128;
				I7x <= 1316;
				I8x <= 857;
				I9x <= 1433;
				I10x <= 1422;
				I11x <= 1762;
				I12x <= 1433;
				I13x <= 1586;
				I14x <= 2068;
				I15x <= 2056;
				I16x <= 2374;
				I17x <= 2221;
				I18x <= 2233;
				I19x <= 2820;
				I20x <= 2938;
				I21x <= 3243;
				I22x <= 3384;
				I23x <= 3232;
				I24x <= 3855;
				I25x <= 3890;
				I26x <= 3960;
				I27x <= 3702;
				I28x <= 3337;
				I29x <= 3678;
				I30x <= 3373;
				I31x <= 3702;
				I32x <= 3349;
				I33x <= 3079;
				I34x <= 3149;
				I35x <= 3208;
				I36x <= 3337;
				I37x <= 3032;
				I38x <= 2538;
				I39x <= 2515;
				I40x <= 2468;
				I41x <= 2421;
				I42x <= 2432;
				I43x <= 2127;
				I44x <= 2409;
				I45x <= 2315;
				I46x <= 2832;
				I47x <= 2538;
				I48x <= 2338;
				I49x <= 2632;
				I50x <= 2233;
				I51x <= 2479;
				I52x <= 2150;
				I53x <= 1962;
				I54x <= 2362;
				I55x <= 2045;
				I56x <= 2479;
				I57x <= 2667;
				I58x <= 2867;
				I59x <= 3902;
				I60x <= 3890;
				I61x <= 3796;
				I62x <= 4572;
				I63x <= 4513;
				I64x <= 4854;
				I65x <= 3196;
				I66x <= 2338;
				I67x <= 1516;
				I68x <= 1210;
				I69x <= 1257;
				I70x <= 669;
				I71x <= 881;
				I72x <= 505;
				I73x <= 658;
				I74x <= 999;
				I75x <= 1057;
				I76x <= 2832;
				I77x <= 5700;
				I78x <= 6699;
				I79x <= 7063;
				I80x <= 7956;
				I81x <= 6840;
				I82x <= 505;
				I83x <= 834;
				I84x <= 1269;
				I85x <= 1093;
				I86x <= 1140;
				I87x <= 987;
				I88x <= 975;
				I89x <= 1210;
				I90x <= 1010;
				I91x <= 1057;
				I92x <= 999;
				I93x <= 893;
				I94x <= 1292;
				I95x <= 1339;
				I96x <= 1539;
				I97x <= 1504;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001100:begin
				I0x <= 8192;
				I1x <= 3512;
				I2x <= 1172;
				I3x <= 87;
				I4x <= 3622;
				I5x <= 4714;
				I6x <= 5085;
				I7x <= 5341;
				I8x <= 5231;
				I9x <= 5370;
				I10x <= 5213;
				I11x <= 5271;
				I12x <= 5527;
				I13x <= 5376;
				I14x <= 5614;
				I15x <= 5503;
				I16x <= 5492;
				I17x <= 5666;
				I18x <= 5492;
				I19x <= 5643;
				I20x <= 5498;
				I21x <= 5561;
				I22x <= 5875;
				I23x <= 5805;
				I24x <= 5950;
				I25x <= 5881;
				I26x <= 5939;
				I27x <= 6334;
				I28x <= 6241;
				I29x <= 6607;
				I30x <= 6577;
				I31x <= 6583;
				I32x <= 6821;
				I33x <= 6607;
				I34x <= 6583;
				I35x <= 6171;
				I36x <= 5869;
				I37x <= 5770;
				I38x <= 5329;
				I39x <= 5347;
				I40x <= 5074;
				I41x <= 4975;
				I42x <= 5074;
				I43x <= 5039;
				I44x <= 5062;
				I45x <= 4952;
				I46x <= 4969;
				I47x <= 5114;
				I48x <= 4871;
				I49x <= 5074;
				I50x <= 4876;
				I51x <= 4963;
				I52x <= 5149;
				I53x <= 5097;
				I54x <= 5196;
				I55x <= 5068;
				I56x <= 5155;
				I57x <= 5242;
				I58x <= 5056;
				I59x <= 5184;
				I60x <= 5027;
				I61x <= 5097;
				I62x <= 5231;
				I63x <= 4975;
				I64x <= 5167;
				I65x <= 5074;
				I66x <= 5149;
				I67x <= 5225;
				I68x <= 5022;
				I69x <= 5056;
				I70x <= 5033;
				I71x <= 5080;
				I72x <= 5190;
				I73x <= 4905;
				I74x <= 4946;
				I75x <= 4853;
				I76x <= 4969;
				I77x <= 5091;
				I78x <= 4905;
				I79x <= 4998;
				I80x <= 4871;
				I81x <= 5016;
				I82x <= 4992;
				I83x <= 4789;
				I84x <= 4975;
				I85x <= 4789;
				I86x <= 4992;
				I87x <= 5091;
				I88x <= 4946;
				I89x <= 5231;
				I90x <= 5416;
				I91x <= 5753;
				I92x <= 5701;
				I93x <= 5800;
				I94x <= 6223;
				I95x <= 5858;
				I96x <= 5649;
				I97x <= 5625;
				I98x <= 4911;
				I99x <= 5010;
				I100x <= 4842;
				I101x <= 4842;
				I102x <= 4789;
				I103x <= 4621;
				I104x <= 4696;
				I105x <= 4592;
				I106x <= 4830;
				I107x <= 4656;
				I108x <= 4493;
				I109x <= 5114;
				I110x <= 4894;
				I111x <= 5219;
				I112x <= 5329;
				I113x <= 6363;
				I114x <= 8006;
				I115x <= 3402;
				I116x <= 865;
				I117x <= 0;
				I118x <= 2873;
				I119x <= 4540;
				I120x <= 4836;
				I121x <= 5074;
				I122x <= 5126;
				I123x <= 4958;
				I124x <= 5114;
				I125x <= 5103;
				I126x <= 5172;
				I127x <= 5300;
				I128x <= 5068;
				I129x <= 5306;
				I130x <= 5184;
				I131x <= 5440;
				I132x <= 5393;
				I133x <= 5213;
				I134x <= 5445;
				I135x <= 5335;
				I136x <= 5567;
				I137x <= 5515;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001101:begin
				I0x <= 8192;
				I1x <= 4262;
				I2x <= 1582;
				I3x <= 0;
				I4x <= 1513;
				I5x <= 1614;
				I6x <= 801;
				I7x <= 1767;
				I8x <= 727;
				I9x <= 1276;
				I10x <= 1434;
				I11x <= 696;
				I12x <= 1751;
				I13x <= 743;
				I14x <= 1450;
				I15x <= 1640;
				I16x <= 933;
				I17x <= 2073;
				I18x <= 1002;
				I19x <= 1735;
				I20x <= 1962;
				I21x <= 1244;
				I22x <= 2357;
				I23x <= 1345;
				I24x <= 2120;
				I25x <= 2299;
				I26x <= 1761;
				I27x <= 2975;
				I28x <= 2073;
				I29x <= 2927;
				I30x <= 3328;
				I31x <= 2669;
				I32x <= 3718;
				I33x <= 2737;
				I34x <= 3265;
				I35x <= 3112;
				I36x <= 2131;
				I37x <= 2806;
				I38x <= 1598;
				I39x <= 2041;
				I40x <= 1935;
				I41x <= 1134;
				I42x <= 2215;
				I43x <= 1128;
				I44x <= 1856;
				I45x <= 1999;
				I46x <= 1329;
				I47x <= 2421;
				I48x <= 1440;
				I49x <= 2141;
				I50x <= 2194;
				I51x <= 1566;
				I52x <= 2626;
				I53x <= 1598;
				I54x <= 2284;
				I55x <= 2284;
				I56x <= 1561;
				I57x <= 2500;
				I58x <= 1476;
				I59x <= 2152;
				I60x <= 2241;
				I61x <= 1450;
				I62x <= 2458;
				I63x <= 1244;
				I64x <= 1909;
				I65x <= 1914;
				I66x <= 1165;
				I67x <= 2210;
				I68x <= 1102;
				I69x <= 1893;
				I70x <= 1898;
				I71x <= 1234;
				I72x <= 2236;
				I73x <= 1086;
				I74x <= 1830;
				I75x <= 1804;
				I76x <= 1134;
				I77x <= 2152;
				I78x <= 1086;
				I79x <= 1909;
				I80x <= 2120;
				I81x <= 1830;
				I82x <= 3011;
				I83x <= 2305;
				I84x <= 3128;
				I85x <= 3402;
				I86x <= 2695;
				I87x <= 3623;
				I88x <= 2452;
				I89x <= 3096;
				I90x <= 2880;
				I91x <= 2004;
				I92x <= 2526;
				I93x <= 1229;
				I94x <= 1809;
				I95x <= 1687;
				I96x <= 996;
				I97x <= 1935;
				I98x <= 875;
				I99x <= 1661;
				I100x <= 1556;
				I101x <= 949;
				I102x <= 1978;
				I103x <= 970;
				I104x <= 1788;
				I105x <= 1756;
				I106x <= 1239;
				I107x <= 2579;
				I108x <= 2458;
				I109x <= 4183;
				I110x <= 6319;
				I111x <= 7859;
				I112x <= 6118;
				I113x <= 1360;
				I114x <= 1461;
				I115x <= 2326;
				I116x <= 1846;
				I117x <= 2632;
				I118x <= 1550;
				I119x <= 2331;
				I120x <= 2215;
				I121x <= 1640;
				I122x <= 2716;
				I123x <= 1709;
				I124x <= 2468;
				I125x <= 2400;
				I126x <= 1904;
				I127x <= 2948;
				I128x <= 1946;
				I129x <= 2853;
				I130x <= 2811;
				I131x <= 2273;
				I132x <= 3317;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001110:begin
				I0x <= 7389;
				I1x <= 5229;
				I2x <= 2555;
				I3x <= 779;
				I4x <= 395;
				I5x <= 443;
				I6x <= 51;
				I7x <= 67;
				I8x <= 90;
				I9x <= 0;
				I10x <= 185;
				I11x <= 229;
				I12x <= 150;
				I13x <= 205;
				I14x <= 122;
				I15x <= 308;
				I16x <= 292;
				I17x <= 320;
				I18x <= 427;
				I19x <= 371;
				I20x <= 458;
				I21x <= 557;
				I22x <= 506;
				I23x <= 609;
				I24x <= 779;
				I25x <= 969;
				I26x <= 1131;
				I27x <= 1281;
				I28x <= 1325;
				I29x <= 1329;
				I30x <= 1467;
				I31x <= 1617;
				I32x <= 1649;
				I33x <= 1574;
				I34x <= 1629;
				I35x <= 1605;
				I36x <= 1507;
				I37x <= 1158;
				I38x <= 1139;
				I39x <= 802;
				I40x <= 700;
				I41x <= 648;
				I42x <= 553;
				I43x <= 371;
				I44x <= 458;
				I45x <= 518;
				I46x <= 581;
				I47x <= 431;
				I48x <= 522;
				I49x <= 411;
				I50x <= 522;
				I51x <= 727;
				I52x <= 494;
				I53x <= 530;
				I54x <= 565;
				I55x <= 632;
				I56x <= 593;
				I57x <= 581;
				I58x <= 514;
				I59x <= 443;
				I60x <= 490;
				I61x <= 597;
				I62x <= 367;
				I63x <= 348;
				I64x <= 403;
				I65x <= 458;
				I66x <= 371;
				I67x <= 423;
				I68x <= 423;
				I69x <= 257;
				I70x <= 312;
				I71x <= 565;
				I72x <= 316;
				I73x <= 324;
				I74x <= 363;
				I75x <= 478;
				I76x <= 688;
				I77x <= 783;
				I78x <= 921;
				I79x <= 945;
				I80x <= 945;
				I81x <= 1427;
				I82x <= 1321;
				I83x <= 1162;
				I84x <= 862;
				I85x <= 609;
				I86x <= 474;
				I87x <= 304;
				I88x <= 158;
				I89x <= 90;
				I90x <= 233;
				I91x <= 249;
				I92x <= 213;
				I93x <= 197;
				I94x <= 193;
				I95x <= 217;
				I96x <= 197;
				I97x <= 75;
				I98x <= 241;
				I99x <= 1186;
				I100x <= 4639;
				I101x <= 8192;
				I102x <= 6499;
				I103x <= 3987;
				I104x <= 1681;
				I105x <= 791;
				I106x <= 715;
				I107x <= 676;
				I108x <= 237;
				I109x <= 213;
				I110x <= 328;
				I111x <= 316;
				I112x <= 356;
				I113x <= 288;
				I114x <= 371;
				I115x <= 292;
				I116x <= 573;
				I117x <= 494;
				I118x <= 403;
				I119x <= 427;
				I120x <= 632;
				I121x <= 751;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01001111:begin
				I0x <= 7598;
				I1x <= 5174;
				I2x <= 2658;
				I3x <= 2048;
				I4x <= 1443;
				I5x <= 855;
				I6x <= 691;
				I7x <= 495;
				I8x <= 462;
				I9x <= 446;
				I10x <= 599;
				I11x <= 691;
				I12x <= 479;
				I13x <= 648;
				I14x <= 697;
				I15x <= 669;
				I16x <= 778;
				I17x <= 936;
				I18x <= 942;
				I19x <= 936;
				I20x <= 1122;
				I21x <= 1154;
				I22x <= 1040;
				I23x <= 1394;
				I24x <= 1465;
				I25x <= 1568;
				I26x <= 1737;
				I27x <= 1988;
				I28x <= 2086;
				I29x <= 2167;
				I30x <= 2097;
				I31x <= 2260;
				I32x <= 2173;
				I33x <= 1939;
				I34x <= 1530;
				I35x <= 1209;
				I36x <= 904;
				I37x <= 757;
				I38x <= 697;
				I39x <= 512;
				I40x <= 675;
				I41x <= 740;
				I42x <= 735;
				I43x <= 424;
				I44x <= 768;
				I45x <= 833;
				I46x <= 964;
				I47x <= 964;
				I48x <= 942;
				I49x <= 860;
				I50x <= 789;
				I51x <= 800;
				I52x <= 795;
				I53x <= 789;
				I54x <= 746;
				I55x <= 653;
				I56x <= 822;
				I57x <= 800;
				I58x <= 648;
				I59x <= 909;
				I60x <= 648;
				I61x <= 626;
				I62x <= 555;
				I63x <= 675;
				I64x <= 626;
				I65x <= 620;
				I66x <= 708;
				I67x <= 561;
				I68x <= 550;
				I69x <= 424;
				I70x <= 484;
				I71x <= 386;
				I72x <= 501;
				I73x <= 364;
				I74x <= 457;
				I75x <= 310;
				I76x <= 326;
				I77x <= 108;
				I78x <= 375;
				I79x <= 386;
				I80x <= 359;
				I81x <= 561;
				I82x <= 708;
				I83x <= 1034;
				I84x <= 991;
				I85x <= 1165;
				I86x <= 1661;
				I87x <= 1595;
				I88x <= 1846;
				I89x <= 1841;
				I90x <= 1230;
				I91x <= 1045;
				I92x <= 686;
				I93x <= 283;
				I94x <= 266;
				I95x <= 81;
				I96x <= 130;
				I97x <= 81;
				I98x <= 157;
				I99x <= 0;
				I100x <= 21;
				I101x <= 185;
				I102x <= 1024;
				I103x <= 3159;
				I104x <= 5196;
				I105x <= 8192;
				I106x <= 5414;
				I107x <= 2598;
				I108x <= 1868;
				I109x <= 1334;
				I110x <= 757;
				I111x <= 326;
				I112x <= 386;
				I113x <= 326;
				I114x <= 261;
				I115x <= 337;
				I116x <= 332;
				I117x <= 315;
				I118x <= 512;
				I119x <= 430;
				I120x <= 577;
				I121x <= 495;
				I122x <= 550;
				I123x <= 735;
				I124x <= 631;
				I125x <= 920;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010000:begin
				I0x <= 8192;
				I1x <= 4079;
				I2x <= 1807;
				I3x <= 835;
				I4x <= 0;
				I5x <= 1310;
				I6x <= 1829;
				I7x <= 2184;
				I8x <= 2162;
				I9x <= 2217;
				I10x <= 2195;
				I11x <= 2146;
				I12x <= 2255;
				I13x <= 2304;
				I14x <= 2381;
				I15x <= 2337;
				I16x <= 2244;
				I17x <= 2217;
				I18x <= 2244;
				I19x <= 2271;
				I20x <= 2266;
				I21x <= 2113;
				I22x <= 2146;
				I23x <= 2118;
				I24x <= 2108;
				I25x <= 2118;
				I26x <= 2086;
				I27x <= 2195;
				I28x <= 2157;
				I29x <= 2293;
				I30x <= 2151;
				I31x <= 2222;
				I32x <= 2282;
				I33x <= 2353;
				I34x <= 2304;
				I35x <= 2512;
				I36x <= 2594;
				I37x <= 2643;
				I38x <= 2626;
				I39x <= 2796;
				I40x <= 2774;
				I41x <= 2883;
				I42x <= 2965;
				I43x <= 2998;
				I44x <= 2905;
				I45x <= 2861;
				I46x <= 2670;
				I47x <= 2566;
				I48x <= 2435;
				I49x <= 2260;
				I50x <= 2408;
				I51x <= 2211;
				I52x <= 2162;
				I53x <= 2118;
				I54x <= 2086;
				I55x <= 2086;
				I56x <= 2037;
				I57x <= 2086;
				I58x <= 2195;
				I59x <= 2135;
				I60x <= 2173;
				I61x <= 2162;
				I62x <= 2195;
				I63x <= 2271;
				I64x <= 2255;
				I65x <= 2255;
				I66x <= 2200;
				I67x <= 2260;
				I68x <= 2184;
				I69x <= 2260;
				I70x <= 2189;
				I71x <= 2075;
				I72x <= 2091;
				I73x <= 2179;
				I74x <= 2233;
				I75x <= 2200;
				I76x <= 2069;
				I77x <= 2108;
				I78x <= 2195;
				I79x <= 2293;
				I80x <= 2288;
				I81x <= 2168;
				I82x <= 2271;
				I83x <= 2250;
				I84x <= 2293;
				I85x <= 2222;
				I86x <= 2179;
				I87x <= 2151;
				I88x <= 2042;
				I89x <= 2053;
				I90x <= 2129;
				I91x <= 2026;
				I92x <= 2157;
				I93x <= 2168;
				I94x <= 2222;
				I95x <= 2222;
				I96x <= 2402;
				I97x <= 2452;
				I98x <= 2632;
				I99x <= 2839;
				I100x <= 3009;
				I101x <= 3402;
				I102x <= 3631;
				I103x <= 3609;
				I104x <= 3549;
				I105x <= 3440;
				I106x <= 3528;
				I107x <= 3129;
				I108x <= 2523;
				I109x <= 2315;
				I110x <= 2058;
				I111x <= 2004;
				I112x <= 1982;
				I113x <= 1927;
				I114x <= 1916;
				I115x <= 1955;
				I116x <= 1884;
				I117x <= 1906;
				I118x <= 2031;
				I119x <= 2424;
				I120x <= 3386;
				I121x <= 4150;
				I122x <= 6662;
				I123x <= 7962;
				I124x <= 3779;
				I125x <= 1856;
				I126x <= 567;
				I127x <= 688;
				I128x <= 1567;
				I129x <= 2042;
				I130x <= 2266;
				I131x <= 2217;
				I132x <= 2353;
				I133x <= 2342;
				I134x <= 2359;
				I135x <= 2342;
				I136x <= 2288;
				I137x <= 2282;
				I138x <= 2271;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010001:begin
				I0x <= 8192;
				I1x <= 6153;
				I2x <= 3917;
				I3x <= 2252;
				I4x <= 0;
				I5x <= 124;
				I6x <= 498;
				I7x <= 1157;
				I8x <= 2419;
				I9x <= 3792;
				I10x <= 4215;
				I11x <= 4350;
				I12x <= 4441;
				I13x <= 4622;
				I14x <= 4628;
				I15x <= 4589;
				I16x <= 4592;
				I17x <= 4631;
				I18x <= 4727;
				I19x <= 4681;
				I20x <= 4674;
				I21x <= 4661;
				I22x <= 4707;
				I23x <= 4704;
				I24x <= 4674;
				I25x <= 4707;
				I26x <= 4776;
				I27x <= 4727;
				I28x <= 4713;
				I29x <= 4648;
				I30x <= 4648;
				I31x <= 4713;
				I32x <= 4700;
				I33x <= 4713;
				I34x <= 4599;
				I35x <= 4674;
				I36x <= 4707;
				I37x <= 4681;
				I38x <= 4713;
				I39x <= 4654;
				I40x <= 4661;
				I41x <= 4661;
				I42x <= 4494;
				I43x <= 4730;
				I44x <= 4651;
				I45x <= 4582;
				I46x <= 4631;
				I47x <= 4612;
				I48x <= 4609;
				I49x <= 4572;
				I50x <= 4448;
				I51x <= 4579;
				I52x <= 4530;
				I53x <= 4566;
				I54x <= 4592;
				I55x <= 4586;
				I56x <= 4622;
				I57x <= 4540;
				I58x <= 4599;
				I59x <= 4586;
				I60x <= 4645;
				I61x <= 4572;
				I62x <= 4609;
				I63x <= 4599;
				I64x <= 4648;
				I65x <= 4599;
				I66x <= 4602;
				I67x <= 4523;
				I68x <= 4599;
				I69x <= 4602;
				I70x <= 4579;
				I71x <= 4520;
				I72x <= 4491;
				I73x <= 4530;
				I74x <= 4523;
				I75x <= 4494;
				I76x <= 4586;
				I77x <= 4484;
				I78x <= 4484;
				I79x <= 4435;
				I80x <= 4530;
				I81x <= 4491;
				I82x <= 4563;
				I83x <= 4402;
				I84x <= 4546;
				I85x <= 4448;
				I86x <= 4441;
				I87x <= 4432;
				I88x <= 4284;
				I89x <= 4497;
				I90x <= 4425;
				I91x <= 4386;
				I92x <= 4497;
				I93x <= 4399;
				I94x <= 4428;
				I95x <= 4379;
				I96x <= 4274;
				I97x <= 4271;
				I98x <= 4418;
				I99x <= 4395;
				I100x <= 4353;
				I101x <= 4366;
				I102x <= 4320;
				I103x <= 4281;
				I104x <= 4317;
				I105x <= 4395;
				I106x <= 4382;
				I107x <= 4277;
				I108x <= 4376;
				I109x <= 4418;
				I110x <= 4415;
				I111x <= 4412;
				I112x <= 4369;
				I113x <= 4373;
				I114x <= 4536;
				I115x <= 4763;
				I116x <= 4956;
				I117x <= 4949;
				I118x <= 4615;
				I119x <= 4831;
				I120x <= 4671;
				I121x <= 4609;
				I122x <= 4550;
				I123x <= 4628;
				I124x <= 4602;
				I125x <= 4474;
				I126x <= 4382;
				I127x <= 4225;
				I128x <= 4199;
				I129x <= 4163;
				I130x <= 4114;
				I131x <= 4294;
				I132x <= 4173;
				I133x <= 4143;
				I134x <= 4271;
				I135x <= 4238;
				I136x <= 4133;
				I137x <= 4225;
				I138x <= 4373;
				I139x <= 4212;
				I140x <= 4779;
				I141x <= 5038;
				I142x <= 5490;
				I143x <= 7123;
				I144x <= 7090;
				I145x <= 5238;
				I146x <= 3651;
				I147x <= 1553;
				I148x <= 262;
				I149x <= 373;
				I150x <= 750;
				I151x <= 1560;
				I152x <= 2730;
				I153x <= 3841;
				I154x <= 4153;
				I155x <= 4238;
				I156x <= 4245;
				I157x <= 4333;
				I158x <= 4389;
				I159x <= 4336;
				I160x <= 4343;
				I161x <= 4451;
				I162x <= 4405;
				I163x <= 4445;
				I164x <= 4556;
				I165x <= 4497;
				I166x <= 4445;
				I167x <= 4399;
				I168x <= 4438;
				I169x <= 4494;
				I170x <= 4464;
				I171x <= 4497;
				I172x <= 4513;
				I173x <= 4435;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010010:begin
				I0x <= 8192;
				I1x <= 6042;
				I2x <= 1926;
				I3x <= 0;
				I4x <= 867;
				I5x <= 2298;
				I6x <= 2951;
				I7x <= 3066;
				I8x <= 3215;
				I9x <= 3339;
				I10x <= 3166;
				I11x <= 3364;
				I12x <= 3480;
				I13x <= 3496;
				I14x <= 3538;
				I15x <= 3471;
				I16x <= 3802;
				I17x <= 3852;
				I18x <= 4182;
				I19x <= 4232;
				I20x <= 4182;
				I21x <= 4439;
				I22x <= 4439;
				I23x <= 4968;
				I24x <= 5323;
				I25x <= 5563;
				I26x <= 5761;
				I27x <= 6075;
				I28x <= 6513;
				I29x <= 6670;
				I30x <= 6976;
				I31x <= 7233;
				I32x <= 7373;
				I33x <= 6993;
				I34x <= 6580;
				I35x <= 5753;
				I36x <= 5282;
				I37x <= 4744;
				I38x <= 4224;
				I39x <= 4058;
				I40x <= 3604;
				I41x <= 3562;
				I42x <= 3389;
				I43x <= 3595;
				I44x <= 3513;
				I45x <= 3232;
				I46x <= 3496;
				I47x <= 3546;
				I48x <= 3529;
				I49x <= 3422;
				I50x <= 3075;
				I51x <= 3521;
				I52x <= 3463;
				I53x <= 3438;
				I54x <= 3488;
				I55x <= 3223;
				I56x <= 3323;
				I57x <= 3372;
				I58x <= 3587;
				I59x <= 3918;
				I60x <= 4199;
				I61x <= 4348;
				I62x <= 4389;
				I63x <= 5042;
				I64x <= 4736;
				I65x <= 4100;
				I66x <= 3678;
				I67x <= 3885;
				I68x <= 3521;
				I69x <= 3504;
				I70x <= 3174;
				I71x <= 2984;
				I72x <= 3066;
				I73x <= 3058;
				I74x <= 3017;
				I75x <= 2860;
				I76x <= 2694;
				I77x <= 2174;
				I78x <= 2116;
				I79x <= 3166;
				I80x <= 5116;
				I81x <= 7613;
				I82x <= 3628;
				I83x <= 2116;
				I84x <= 41;
				I85x <= 661;
				I86x <= 2074;
				I87x <= 2777;
				I88x <= 2818;
				I89x <= 3124;
				I90x <= 3199;
				I91x <= 2926;
				I92x <= 3182;
				I93x <= 3207;
				I94x <= 3414;
				I95x <= 3422;
				I96x <= 3496;
				I97x <= 3653;
				I98x <= 3819;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010011:begin
				I0x <= 8192;
				I1x <= 6978;
				I2x <= 3800;
				I3x <= 2934;
				I4x <= 2228;
				I5x <= 2064;
				I6x <= 2198;
				I7x <= 2098;
				I8x <= 2069;
				I9x <= 2049;
				I10x <= 1924;
				I11x <= 2278;
				I12x <= 2347;
				I13x <= 2382;
				I14x <= 2447;
				I15x <= 2392;
				I16x <= 2382;
				I17x <= 2476;
				I18x <= 2342;
				I19x <= 2342;
				I20x <= 2377;
				I21x <= 2442;
				I22x <= 2476;
				I23x <= 2352;
				I24x <= 2442;
				I25x <= 2307;
				I26x <= 2278;
				I27x <= 2138;
				I28x <= 1989;
				I29x <= 2069;
				I30x <= 1949;
				I31x <= 2044;
				I32x <= 1929;
				I33x <= 1999;
				I34x <= 2208;
				I35x <= 2168;
				I36x <= 2287;
				I37x <= 2367;
				I38x <= 2506;
				I39x <= 2641;
				I40x <= 2551;
				I41x <= 2705;
				I42x <= 2760;
				I43x <= 2651;
				I44x <= 2745;
				I45x <= 2755;
				I46x <= 2795;
				I47x <= 2775;
				I48x <= 2740;
				I49x <= 2815;
				I50x <= 2760;
				I51x <= 2755;
				I52x <= 2725;
				I53x <= 2626;
				I54x <= 2675;
				I55x <= 2422;
				I56x <= 2695;
				I57x <= 2715;
				I58x <= 2566;
				I59x <= 2760;
				I60x <= 2601;
				I61x <= 2601;
				I62x <= 2611;
				I63x <= 2666;
				I64x <= 2989;
				I65x <= 3063;
				I66x <= 3466;
				I67x <= 3874;
				I68x <= 3814;
				I69x <= 3685;
				I70x <= 3312;
				I71x <= 3223;
				I72x <= 2755;
				I73x <= 2611;
				I74x <= 2516;
				I75x <= 2268;
				I76x <= 2292;
				I77x <= 2228;
				I78x <= 2143;
				I79x <= 1502;
				I80x <= 0;
				I81x <= 860;
				I82x <= 4541;
				I83x <= 7629;
				I84x <= 8042;
				I85x <= 5754;
				I86x <= 3745;
				I87x <= 2775;
				I88x <= 2292;
				I89x <= 2402;
				I90x <= 2357;
				I91x <= 2382;
				I92x <= 2392;
				I93x <= 2317;
				I94x <= 2506;
				I95x <= 2402;
				I96x <= 2576;
				I97x <= 2616;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010100:begin
				I0x <= 8192;
				I1x <= 3642;
				I2x <= 593;
				I3x <= 508;
				I4x <= 1234;
				I5x <= 1163;
				I6x <= 1057;
				I7x <= 876;
				I8x <= 739;
				I9x <= 863;
				I10x <= 588;
				I11x <= 668;
				I12x <= 827;
				I13x <= 871;
				I14x <= 730;
				I15x <= 663;
				I16x <= 752;
				I17x <= 876;
				I18x <= 655;
				I19x <= 836;
				I20x <= 712;
				I21x <= 876;
				I22x <= 1411;
				I23x <= 947;
				I24x <= 1243;
				I25x <= 1230;
				I26x <= 1575;
				I27x <= 1305;
				I28x <= 1779;
				I29x <= 1779;
				I30x <= 1978;
				I31x <= 2164;
				I32x <= 2234;
				I33x <= 2655;
				I34x <= 2487;
				I35x <= 2416;
				I36x <= 2350;
				I37x <= 2345;
				I38x <= 2177;
				I39x <= 1916;
				I40x <= 1526;
				I41x <= 1402;
				I42x <= 1168;
				I43x <= 1035;
				I44x <= 1146;
				I45x <= 1305;
				I46x <= 606;
				I47x <= 783;
				I48x <= 690;
				I49x <= 619;
				I50x <= 646;
				I51x <= 566;
				I52x <= 694;
				I53x <= 867;
				I54x <= 615;
				I55x <= 893;
				I56x <= 809;
				I57x <= 964;
				I58x <= 752;
				I59x <= 739;
				I60x <= 916;
				I61x <= 951;
				I62x <= 650;
				I63x <= 358;
				I64x <= 522;
				I65x <= 451;
				I66x <= 646;
				I67x <= 460;
				I68x <= 624;
				I69x <= 460;
				I70x <= 677;
				I71x <= 345;
				I72x <= 681;
				I73x <= 893;
				I74x <= 482;
				I75x <= 677;
				I76x <= 1615;
				I77x <= 1248;
				I78x <= 1482;
				I79x <= 1845;
				I80x <= 1464;
				I81x <= 1730;
				I82x <= 1686;
				I83x <= 1394;
				I84x <= 1438;
				I85x <= 991;
				I86x <= 712;
				I87x <= 557;
				I88x <= 0;
				I89x <= 902;
				I90x <= 677;
				I91x <= 641;
				I92x <= 469;
				I93x <= 420;
				I94x <= 544;
				I95x <= 296;
				I96x <= 230;
				I97x <= 544;
				I98x <= 1557;
				I99x <= 4779;
				I100x <= 7359;
				I101x <= 6253;
				I102x <= 1885;
				I103x <= 13;
				I104x <= 491;
				I105x <= 814;
				I106x <= 774;
				I107x <= 544;
				I108x <= 743;
				I109x <= 508;
				I110x <= 575;
				I111x <= 716;
				I112x <= 1026;
				I113x <= 969;
				I114x <= 907;
				I115x <= 893;
				I116x <= 809;
				I117x <= 1256;
				I118x <= 1040;
				I119x <= 1048;
				I120x <= 1053;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010101:begin
				I0x <= 8192;
				I1x <= 3448;
				I2x <= 2989;
				I3x <= 1231;
				I4x <= 1149;
				I5x <= 1265;
				I6x <= 1270;
				I7x <= 1154;
				I8x <= 1149;
				I9x <= 1207;
				I10x <= 1231;
				I11x <= 1251;
				I12x <= 1313;
				I13x <= 1308;
				I14x <= 1347;
				I15x <= 1381;
				I16x <= 1434;
				I17x <= 1516;
				I18x <= 1516;
				I19x <= 1492;
				I20x <= 1627;
				I21x <= 1719;
				I22x <= 1700;
				I23x <= 1830;
				I24x <= 1888;
				I25x <= 2043;
				I26x <= 2159;
				I27x <= 2221;
				I28x <= 2279;
				I29x <= 2241;
				I30x <= 2159;
				I31x <= 1990;
				I32x <= 1859;
				I33x <= 1637;
				I34x <= 1482;
				I35x <= 1400;
				I36x <= 1270;
				I37x <= 1231;
				I38x <= 1222;
				I39x <= 1154;
				I40x <= 1222;
				I41x <= 1173;
				I42x <= 1207;
				I43x <= 1226;
				I44x <= 1275;
				I45x <= 1289;
				I46x <= 1352;
				I47x <= 1371;
				I48x <= 1424;
				I49x <= 1458;
				I50x <= 1415;
				I51x <= 1362;
				I52x <= 1323;
				I53x <= 1313;
				I54x <= 1318;
				I55x <= 1299;
				I56x <= 1328;
				I57x <= 1294;
				I58x <= 1299;
				I59x <= 1318;
				I60x <= 1280;
				I61x <= 1337;
				I62x <= 1598;
				I63x <= 1912;
				I64x <= 1956;
				I65x <= 2076;
				I66x <= 1990;
				I67x <= 2091;
				I68x <= 1598;
				I69x <= 1632;
				I70x <= 1236;
				I71x <= 1115;
				I72x <= 1139;
				I73x <= 995;
				I74x <= 883;
				I75x <= 825;
				I76x <= 912;
				I77x <= 864;
				I78x <= 507;
				I79x <= 0;
				I80x <= 1743;
				I81x <= 6134;
				I82x <= 7230;
				I83x <= 3361;
				I84x <= 2052;
				I85x <= 1120;
				I86x <= 1043;
				I87x <= 1231;
				I88x <= 1062;
				I89x <= 1135;
				I90x <= 1183;
				I91x <= 1164;
				I92x <= 1096;
				I93x <= 1130;
				I94x <= 1236;
				I95x <= 1202;
				I96x <= 1313;
				I97x <= 1260;
				I98x <= 1294;
				I99x <= 1342;
				I100x <= 1400;
				I101x <= 1627;
				I102x <= 1584;
				I103x <= 1647;
				I104x <= 1825;
				I105x <= 1801;
				I106x <= 1912;
				I107x <= 1922;
				I108x <= 1985;
				I109x <= 2101;
				I110x <= 2168;
				I111x <= 2120;
				I112x <= 1980;
				I113x <= 1883;
				I114x <= 1685;
				I115x <= 1540;
				I116x <= 1381;
				I117x <= 1226;
				I118x <= 1197;
				I119x <= 1130;
				I120x <= 1188;
				I121x <= 1226;
				I122x <= 1231;
				I123x <= 1154;
				I124x <= 1154;
				I125x <= 1110;
				I126x <= 1222;
				I127x <= 1328;
				I128x <= 1241;
				I129x <= 1308;
				I130x <= 1251;
				I131x <= 1280;
				I132x <= 1280;
				I133x <= 1318;
				I134x <= 1318;
				I135x <= 1212;
				I136x <= 1231;
				I137x <= 1236;
				I138x <= 1207;
				I139x <= 1120;
				I140x <= 1183;
				I141x <= 1197;
				I142x <= 1154;
				I143x <= 1299;
				I144x <= 1690;
				I145x <= 1714;
				I146x <= 1912;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010110:begin
				I0x <= 8192;
				I1x <= 5736;
				I2x <= 1112;
				I3x <= 828;
				I4x <= 1116;
				I5x <= 1198;
				I6x <= 1177;
				I7x <= 1221;
				I8x <= 1179;
				I9x <= 1189;
				I10x <= 1123;
				I11x <= 1096;
				I12x <= 1006;
				I13x <= 1045;
				I14x <= 1068;
				I15x <= 1016;
				I16x <= 991;
				I17x <= 1027;
				I18x <= 1085;
				I19x <= 1083;
				I20x <= 1091;
				I21x <= 1123;
				I22x <= 1146;
				I23x <= 1329;
				I24x <= 1369;
				I25x <= 1413;
				I26x <= 1599;
				I27x <= 1626;
				I28x <= 1784;
				I29x <= 1770;
				I30x <= 1816;
				I31x <= 1820;
				I32x <= 1880;
				I33x <= 1943;
				I34x <= 1901;
				I35x <= 1891;
				I36x <= 1910;
				I37x <= 1801;
				I38x <= 1839;
				I39x <= 1849;
				I40x <= 1778;
				I41x <= 1789;
				I42x <= 1730;
				I43x <= 1772;
				I44x <= 1755;
				I45x <= 1724;
				I46x <= 1722;
				I47x <= 1649;
				I48x <= 1638;
				I49x <= 1651;
				I50x <= 1553;
				I51x <= 1580;
				I52x <= 1588;
				I53x <= 1557;
				I54x <= 1546;
				I55x <= 1538;
				I56x <= 1567;
				I57x <= 1501;
				I58x <= 1553;
				I59x <= 1657;
				I60x <= 1853;
				I61x <= 1972;
				I62x <= 1999;
				I63x <= 2018;
				I64x <= 1943;
				I65x <= 1914;
				I66x <= 1855;
				I67x <= 1684;
				I68x <= 1607;
				I69x <= 1532;
				I70x <= 1384;
				I71x <= 1601;
				I72x <= 1411;
				I73x <= 1455;
				I74x <= 1453;
				I75x <= 1421;
				I76x <= 1444;
				I77x <= 1409;
				I78x <= 1492;
				I79x <= 1430;
				I80x <= 1064;
				I81x <= 659;
				I82x <= 0;
				I83x <= 878;
				I84x <= 4068;
				I85x <= 7956;
				I86x <= 4870;
				I87x <= 918;
				I88x <= 659;
				I89x <= 914;
				I90x <= 947;
				I91x <= 1016;
				I92x <= 943;
				I93x <= 1027;
				I94x <= 1006;
				I95x <= 916;
				I96x <= 974;
				I97x <= 868;
				I98x <= 901;
				I99x <= 910;
				I100x <= 835;
				I101x <= 851;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01010111:begin
				I0x <= 8192;
				I1x <= 6411;
				I2x <= 4661;
				I3x <= 3676;
				I4x <= 3236;
				I5x <= 2671;
				I6x <= 2545;
				I7x <= 2702;
				I8x <= 2964;
				I9x <= 2618;
				I10x <= 2985;
				I11x <= 2629;
				I12x <= 3037;
				I13x <= 2755;
				I14x <= 2817;
				I15x <= 3184;
				I16x <= 2681;
				I17x <= 3017;
				I18x <= 3079;
				I19x <= 2859;
				I20x <= 3048;
				I21x <= 2859;
				I22x <= 2828;
				I23x <= 2943;
				I24x <= 2912;
				I25x <= 2755;
				I26x <= 2199;
				I27x <= 2304;
				I28x <= 1906;
				I29x <= 1361;
				I30x <= 1120;
				I31x <= 597;
				I32x <= 576;
				I33x <= 0;
				I34x <= 41;
				I35x <= 199;
				I36x <= 0;
				I37x <= 639;
				I38x <= 628;
				I39x <= 806;
				I40x <= 921;
				I41x <= 775;
				I42x <= 1047;
				I43x <= 1005;
				I44x <= 1215;
				I45x <= 1099;
				I46x <= 722;
				I47x <= 1005;
				I48x <= 817;
				I49x <= 879;
				I50x <= 911;
				I51x <= 670;
				I52x <= 838;
				I53x <= 733;
				I54x <= 743;
				I55x <= 523;
				I56x <= 240;
				I57x <= 911;
				I58x <= 628;
				I59x <= 0;
				I60x <= 0;
				I61x <= 0;
				I62x <= 0;
				I63x <= 0;
				I64x <= 0;
				I65x <= 0;
				I66x <= 0;
				I67x <= 0;
				I68x <= 0;
				I69x <= 0;
				I70x <= 0;
				I71x <= 0;
				I72x <= 0;
				I73x <= 0;
				I74x <= 0;
				I75x <= 0;
				I76x <= 0;
				I77x <= 0;
				I78x <= 0;
				I79x <= 0;
				I80x <= 0;
				I81x <= 0;
				I82x <= 0;
				I83x <= 0;
				I84x <= 0;
				I85x <= 0;
				I86x <= 0;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011000:begin
				I0x <= 8192;
				I1x <= 2922;
				I2x <= 1968;
				I3x <= 2078;
				I4x <= 85;
				I5x <= 293;
				I6x <= 0;
				I7x <= 660;
				I8x <= 452;
				I9x <= 550;
				I10x <= 672;
				I11x <= 281;
				I12x <= 513;
				I13x <= 403;
				I14x <= 537;
				I15x <= 623;
				I16x <= 684;
				I17x <= 1369;
				I18x <= 1222;
				I19x <= 1357;
				I20x <= 1601;
				I21x <= 1528;
				I22x <= 2115;
				I23x <= 1956;
				I24x <= 2310;
				I25x <= 2579;
				I26x <= 2494;
				I27x <= 3044;
				I28x <= 2799;
				I29x <= 2799;
				I30x <= 2677;
				I31x <= 2151;
				I32x <= 2274;
				I33x <= 1687;
				I34x <= 1491;
				I35x <= 1675;
				I36x <= 1283;
				I37x <= 1503;
				I38x <= 1222;
				I39x <= 1357;
				I40x <= 1540;
				I41x <= 1308;
				I42x <= 1748;
				I43x <= 1589;
				I44x <= 1613;
				I45x <= 1980;
				I46x <= 1785;
				I47x <= 2347;
				I48x <= 2041;
				I49x <= 2029;
				I50x <= 2188;
				I51x <= 1723;
				I52x <= 2078;
				I53x <= 1626;
				I54x <= 1821;
				I55x <= 1748;
				I56x <= 1393;
				I57x <= 1809;
				I58x <= 1540;
				I59x <= 1662;
				I60x <= 1723;
				I61x <= 1393;
				I62x <= 2543;
				I63x <= 3081;
				I64x <= 3533;
				I65x <= 3912;
				I66x <= 4181;
				I67x <= 4902;
				I68x <= 4010;
				I69x <= 4572;
				I70x <= 4866;
				I71x <= 4169;
				I72x <= 3558;
				I73x <= 1821;
				I74x <= 1198;
				I75x <= 1283;
				I76x <= 880;
				I77x <= 1088;
				I78x <= 574;
				I79x <= 1748;
				I80x <= 1418;
				I81x <= 452;
				I82x <= 3484;
				I83x <= 7996;
				I84x <= 4377;
				I85x <= 2457;
				I86x <= 2983;
				I87x <= 917;
				I88x <= 599;
				I89x <= 623;
				I90x <= 904;
				I91x <= 990;
				I92x <= 1442;
				I93x <= 1051;
				I94x <= 1075;
				I95x <= 1393;
				I96x <= 1112;
				I97x <= 1491;
				I98x <= 1283;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011001:begin
				I0x <= 7672;
				I1x <= 7623;
				I2x <= 4370;
				I3x <= 1587;
				I4x <= 2092;
				I5x <= 1464;
				I6x <= 867;
				I7x <= 930;
				I8x <= 1019;
				I9x <= 1156;
				I10x <= 1121;
				I11x <= 1337;
				I12x <= 1298;
				I13x <= 1460;
				I14x <= 1714;
				I15x <= 1724;
				I16x <= 2234;
				I17x <= 1896;
				I18x <= 2013;
				I19x <= 2302;
				I20x <= 1994;
				I21x <= 2278;
				I22x <= 2033;
				I23x <= 1852;
				I24x <= 1984;
				I25x <= 1607;
				I26x <= 1827;
				I27x <= 1729;
				I28x <= 1685;
				I29x <= 2033;
				I30x <= 1626;
				I31x <= 1935;
				I32x <= 1964;
				I33x <= 1832;
				I34x <= 2052;
				I35x <= 1788;
				I36x <= 2082;
				I37x <= 1705;
				I38x <= 1807;
				I39x <= 1852;
				I40x <= 1509;
				I41x <= 1773;
				I42x <= 1641;
				I43x <= 1553;
				I44x <= 1719;
				I45x <= 2082;
				I46x <= 2537;
				I47x <= 2557;
				I48x <= 2724;
				I49x <= 2778;
				I50x <= 2322;
				I51x <= 2400;
				I52x <= 1950;
				I53x <= 1935;
				I54x <= 2082;
				I55x <= 1950;
				I56x <= 1602;
				I57x <= 1381;
				I58x <= 1332;
				I59x <= 1411;
				I60x <= 1161;
				I61x <= 1450;
				I62x <= 1268;
				I63x <= 681;
				I64x <= 916;
				I65x <= 0;
				I66x <= 480;
				I67x <= 3522;
				I68x <= 7731;
				I69x <= 8192;
				I70x <= 4840;
				I71x <= 2082;
				I72x <= 2302;
				I73x <= 2302;
				I74x <= 1406;
				I75x <= 1489;
				I76x <= 1852;
				I77x <= 1401;
				I78x <= 1847;
				I79x <= 1876;
				I80x <= 1783;
				I81x <= 0;
				I82x <= 0;
				I83x <= 0;
				I84x <= 0;
				I85x <= 0;
				I86x <= 0;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011010:begin
				I0x <= 7955;
				I1x <= 4858;
				I2x <= 1278;
				I3x <= 0;
				I4x <= 191;
				I5x <= 881;
				I6x <= 2371;
				I7x <= 2829;
				I8x <= 2789;
				I9x <= 2940;
				I10x <= 3031;
				I11x <= 3041;
				I12x <= 3252;
				I13x <= 3388;
				I14x <= 3454;
				I15x <= 3454;
				I16x <= 3564;
				I17x <= 3786;
				I18x <= 3569;
				I19x <= 3806;
				I20x <= 3851;
				I21x <= 3836;
				I22x <= 3982;
				I23x <= 4038;
				I24x <= 4063;
				I25x <= 3937;
				I26x <= 3801;
				I27x <= 3861;
				I28x <= 3776;
				I29x <= 3625;
				I30x <= 3519;
				I31x <= 3277;
				I32x <= 3257;
				I33x <= 3222;
				I34x <= 3212;
				I35x <= 3167;
				I36x <= 3106;
				I37x <= 3031;
				I38x <= 3146;
				I39x <= 3131;
				I40x <= 3242;
				I41x <= 3212;
				I42x <= 3328;
				I43x <= 3136;
				I44x <= 3398;
				I45x <= 3121;
				I46x <= 3187;
				I47x <= 3338;
				I48x <= 2809;
				I49x <= 3207;
				I50x <= 3242;
				I51x <= 3272;
				I52x <= 3423;
				I53x <= 3257;
				I54x <= 3308;
				I55x <= 3469;
				I56x <= 3408;
				I57x <= 3529;
				I58x <= 3187;
				I59x <= 3564;
				I60x <= 3438;
				I61x <= 3343;
				I62x <= 3589;
				I63x <= 3549;
				I64x <= 4083;
				I65x <= 4340;
				I66x <= 4491;
				I67x <= 4732;
				I68x <= 5019;
				I69x <= 5009;
				I70x <= 4959;
				I71x <= 4345;
				I72x <= 4395;
				I73x <= 4365;
				I74x <= 4294;
				I75x <= 3947;
				I76x <= 3287;
				I77x <= 3509;
				I78x <= 3398;
				I79x <= 3438;
				I80x <= 3358;
				I81x <= 3272;
				I82x <= 3589;
				I83x <= 2910;
				I84x <= 4204;
				I85x <= 8192;
				I86x <= 6605;
				I87x <= 2789;
				I88x <= 251;
				I89x <= 518;
				I90x <= 805;
				I91x <= 2895;
				I92x <= 3489;
				I93x <= 3584;
				I94x <= 3922;
				I95x <= 3600;
				I96x <= 3861;
				I97x <= 3957;
				I98x <= 3892;
				I99x <= 3957;
				I100x <= 4043;
				I101x <= 4063;
				I102x <= 4340;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011011:begin
				I0x <= 8192;
				I1x <= 5302;
				I2x <= 470;
				I3x <= 1360;
				I4x <= 1610;
				I5x <= 1022;
				I6x <= 941;
				I7x <= 933;
				I8x <= 860;
				I9x <= 853;
				I10x <= 1066;
				I11x <= 1051;
				I12x <= 992;
				I13x <= 1051;
				I14x <= 1095;
				I15x <= 1110;
				I16x <= 1132;
				I17x <= 1301;
				I18x <= 1242;
				I19x <= 1588;
				I20x <= 1610;
				I21x <= 1588;
				I22x <= 1706;
				I23x <= 1654;
				I24x <= 1632;
				I25x <= 1757;
				I26x <= 1889;
				I27x <= 2139;
				I28x <= 2206;
				I29x <= 2301;
				I30x <= 2507;
				I31x <= 2529;
				I32x <= 2566;
				I33x <= 2316;
				I34x <= 2051;
				I35x <= 2051;
				I36x <= 2000;
				I37x <= 1963;
				I38x <= 1639;
				I39x <= 1603;
				I40x <= 1639;
				I41x <= 1875;
				I42x <= 1735;
				I43x <= 1558;
				I44x <= 1507;
				I45x <= 1809;
				I46x <= 1809;
				I47x <= 1581;
				I48x <= 1698;
				I49x <= 1720;
				I50x <= 1691;
				I51x <= 1448;
				I52x <= 1632;
				I53x <= 1691;
				I54x <= 1647;
				I55x <= 1706;
				I56x <= 1676;
				I57x <= 1706;
				I58x <= 1654;
				I59x <= 1529;
				I60x <= 2198;
				I61x <= 2426;
				I62x <= 2992;
				I63x <= 3257;
				I64x <= 3551;
				I65x <= 3456;
				I66x <= 3515;
				I67x <= 3551;
				I68x <= 2654;
				I69x <= 2441;
				I70x <= 2478;
				I71x <= 1963;
				I72x <= 1558;
				I73x <= 1456;
				I74x <= 1367;
				I75x <= 1345;
				I76x <= 1139;
				I77x <= 1198;
				I78x <= 1198;
				I79x <= 1051;
				I80x <= 1654;
				I81x <= 3478;
				I82x <= 5412;
				I83x <= 6221;
				I84x <= 7839;
				I85x <= 5037;
				I86x <= 0;
				I87x <= 1264;
				I88x <= 1632;
				I89x <= 1404;
				I90x <= 1279;
				I91x <= 1183;
				I92x <= 1375;
				I93x <= 1073;
				I94x <= 1206;
				I95x <= 1257;
				I96x <= 1529;
				I97x <= 1573;
				I98x <= 1404;
				I99x <= 1250;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011100:begin
				I0x <= 8192;
				I1x <= 6107;
				I2x <= 2368;
				I3x <= 0;
				I4x <= 1110;
				I5x <= 1687;
				I6x <= 2119;
				I7x <= 3055;
				I8x <= 3528;
				I9x <= 3744;
				I10x <= 3864;
				I11x <= 3908;
				I12x <= 3832;
				I13x <= 3837;
				I14x <= 3845;
				I15x <= 3818;
				I16x <= 3801;
				I17x <= 3788;
				I18x <= 3875;
				I19x <= 3968;
				I20x <= 3982;
				I21x <= 3987;
				I22x <= 4037;
				I23x <= 4171;
				I24x <= 4212;
				I25x <= 4214;
				I26x <= 4351;
				I27x <= 4351;
				I28x <= 4485;
				I29x <= 4425;
				I30x <= 4280;
				I31x <= 4152;
				I32x <= 4132;
				I33x <= 4083;
				I34x <= 4064;
				I35x <= 4004;
				I36x <= 3957;
				I37x <= 3985;
				I38x <= 3974;
				I39x <= 3933;
				I40x <= 3908;
				I41x <= 3897;
				I42x <= 3892;
				I43x <= 3815;
				I44x <= 3837;
				I45x <= 3840;
				I46x <= 3955;
				I47x <= 4100;
				I48x <= 4234;
				I49x <= 4250;
				I50x <= 4307;
				I51x <= 4307;
				I52x <= 4165;
				I53x <= 4050;
				I54x <= 3977;
				I55x <= 4018;
				I56x <= 4007;
				I57x <= 3927;
				I58x <= 3916;
				I59x <= 3960;
				I60x <= 4059;
				I61x <= 3982;
				I62x <= 4091;
				I63x <= 4064;
				I64x <= 4094;
				I65x <= 4031;
				I66x <= 4455;
				I67x <= 5836;
				I68x <= 6446;
				I69x <= 6118;
				I70x <= 8142;
				I71x <= 6233;
				I72x <= 2636;
				I73x <= 306;
				I74x <= 1299;
				I75x <= 1827;
				I76x <= 2286;
				I77x <= 3077;
				I78x <= 3607;
				I79x <= 3774;
				I80x <= 3941;
				I81x <= 3922;
				I82x <= 3853;
				I83x <= 3812;
				I84x <= 0;
				I85x <= 0;
				I86x <= 0;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011101:begin
				I0x <= 8192;
				I1x <= 5196;
				I2x <= 1563;
				I3x <= 124;
				I4x <= 546;
				I5x <= 1522;
				I6x <= 1722;
				I7x <= 1653;
				I8x <= 1570;
				I9x <= 1812;
				I10x <= 1951;
				I11x <= 2027;
				I12x <= 1978;
				I13x <= 1819;
				I14x <= 2117;
				I15x <= 2158;
				I16x <= 2241;
				I17x <= 2165;
				I18x <= 2117;
				I19x <= 2331;
				I20x <= 2338;
				I21x <= 2449;
				I22x <= 2324;
				I23x <= 2193;
				I24x <= 2546;
				I25x <= 2283;
				I26x <= 2262;
				I27x <= 2068;
				I28x <= 1937;
				I29x <= 2124;
				I30x <= 1930;
				I31x <= 1971;
				I32x <= 1778;
				I33x <= 1577;
				I34x <= 1702;
				I35x <= 1501;
				I36x <= 1494;
				I37x <= 1314;
				I38x <= 1134;
				I39x <= 1439;
				I40x <= 1335;
				I41x <= 1404;
				I42x <= 1300;
				I43x <= 1245;
				I44x <= 1536;
				I45x <= 1425;
				I46x <= 1494;
				I47x <= 1321;
				I48x <= 1231;
				I49x <= 1549;
				I50x <= 1508;
				I51x <= 1964;
				I52x <= 1819;
				I53x <= 1854;
				I54x <= 2511;
				I55x <= 2947;
				I56x <= 3134;
				I57x <= 3175;
				I58x <= 3002;
				I59x <= 3044;
				I60x <= 2220;
				I61x <= 1639;
				I62x <= 1293;
				I63x <= 1093;
				I64x <= 1134;
				I65x <= 899;
				I66x <= 1017;
				I67x <= 906;
				I68x <= 671;
				I69x <= 1646;
				I70x <= 1280;
				I71x <= 1030;
				I72x <= 1349;
				I73x <= 5320;
				I74x <= 5742;
				I75x <= 1632;
				I76x <= 83;
				I77x <= 0;
				I78x <= 726;
				I79x <= 1259;
				I80x <= 1065;
				I81x <= 1286;
				I82x <= 1307;
				I83x <= 1210;
				I84x <= 1542;
				I85x <= 1335;
				I86x <= 1605;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011110:begin
				I0x <= 7568;
				I1x <= 7310;
				I2x <= 6369;
				I3x <= 6090;
				I4x <= 3896;
				I5x <= 1291;
				I6x <= 853;
				I7x <= 0;
				I8x <= 629;
				I9x <= 1346;
				I10x <= 1389;
				I11x <= 1264;
				I12x <= 1121;
				I13x <= 1313;
				I14x <= 1220;
				I15x <= 1236;
				I16x <= 1247;
				I17x <= 1400;
				I18x <= 1253;
				I19x <= 1225;
				I20x <= 1105;
				I21x <= 1127;
				I22x <= 1176;
				I23x <= 1088;
				I24x <= 1187;
				I25x <= 1121;
				I26x <= 1307;
				I27x <= 1099;
				I28x <= 1269;
				I29x <= 1384;
				I30x <= 1258;
				I31x <= 1422;
				I32x <= 1225;
				I33x <= 1220;
				I34x <= 1028;
				I35x <= 612;
				I36x <= 733;
				I37x <= 640;
				I38x <= 738;
				I39x <= 826;
				I40x <= 979;
				I41x <= 1028;
				I42x <= 946;
				I43x <= 1127;
				I44x <= 1488;
				I45x <= 1482;
				I46x <= 1395;
				I47x <= 1597;
				I48x <= 1931;
				I49x <= 1816;
				I50x <= 1909;
				I51x <= 2008;
				I52x <= 2068;
				I53x <= 1849;
				I54x <= 1980;
				I55x <= 2084;
				I56x <= 1898;
				I57x <= 1948;
				I58x <= 1805;
				I59x <= 1948;
				I60x <= 1975;
				I61x <= 1833;
				I62x <= 1964;
				I63x <= 1959;
				I64x <= 2249;
				I65x <= 1849;
				I66x <= 1871;
				I67x <= 2041;
				I68x <= 2008;
				I69x <= 1849;
				I70x <= 1876;
				I71x <= 2057;
				I72x <= 1915;
				I73x <= 2013;
				I74x <= 2095;
				I75x <= 2150;
				I76x <= 2139;
				I77x <= 2249;
				I78x <= 2281;
				I79x <= 2364;
				I80x <= 2489;
				I81x <= 2774;
				I82x <= 2566;
				I83x <= 2451;
				I84x <= 3091;
				I85x <= 2889;
				I86x <= 2659;
				I87x <= 2747;
				I88x <= 2648;
				I89x <= 2637;
				I90x <= 2188;
				I91x <= 2123;
				I92x <= 1986;
				I93x <= 2019;
				I94x <= 2052;
				I95x <= 1959;
				I96x <= 2101;
				I97x <= 2035;
				I98x <= 2457;
				I99x <= 3365;
				I100x <= 5302;
				I101x <= 6506;
				I102x <= 7048;
				I103x <= 8192;
				I104x <= 7261;
				I105x <= 6714;
				I106x <= 5329;
				I107x <= 3130;
				I108x <= 1461;
				I109x <= 788;
				I110x <= 344;
				I111x <= 1444;
				I112x <= 1866;
				I113x <= 1915;
				I114x <= 2079;
				I115x <= 2199;
				I116x <= 2095;
				I117x <= 2134;
				I118x <= 2210;
				I119x <= 2052;
				I120x <= 2095;
				I121x <= 2090;
				I122x <= 2052;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01011111:begin
				I0x <= 8192;
				I1x <= 6685;
				I2x <= 4599;
				I3x <= 3528;
				I4x <= 3084;
				I5x <= 1966;
				I6x <= 2394;
				I7x <= 1102;
				I8x <= 1839;
				I9x <= 1506;
				I10x <= 1181;
				I11x <= 1808;
				I12x <= 1649;
				I13x <= 1927;
				I14x <= 2180;
				I15x <= 1633;
				I16x <= 2283;
				I17x <= 1609;
				I18x <= 2204;
				I19x <= 2410;
				I20x <= 2038;
				I21x <= 2950;
				I22x <= 1705;
				I23x <= 2609;
				I24x <= 2902;
				I25x <= 2038;
				I26x <= 3251;
				I27x <= 2513;
				I28x <= 2656;
				I29x <= 3195;
				I30x <= 2339;
				I31x <= 2799;
				I32x <= 1697;
				I33x <= 2482;
				I34x <= 2228;
				I35x <= 1649;
				I36x <= 2442;
				I37x <= 1292;
				I38x <= 1919;
				I39x <= 2371;
				I40x <= 1649;
				I41x <= 2196;
				I42x <= 1633;
				I43x <= 1847;
				I44x <= 2164;
				I45x <= 1816;
				I46x <= 2513;
				I47x <= 1197;
				I48x <= 1641;
				I49x <= 2220;
				I50x <= 2252;
				I51x <= 3203;
				I52x <= 2418;
				I53x <= 2958;
				I54x <= 3164;
				I55x <= 2474;
				I56x <= 3243;
				I57x <= 1601;
				I58x <= 2053;
				I59x <= 1998;
				I60x <= 1078;
				I61x <= 1705;
				I62x <= 158;
				I63x <= 1126;
				I64x <= 1062;
				I65x <= 499;
				I66x <= 1395;
				I67x <= 333;
				I68x <= 1578;
				I69x <= 1665;
				I70x <= 2180;
				I71x <= 5360;
				I72x <= 8112;
				I73x <= 5313;
				I74x <= 4131;
				I75x <= 2910;
				I76x <= 2965;
				I77x <= 1340;
				I78x <= 1546;
				I79x <= 1023;
				I80x <= 0;
				I81x <= 1252;
				I82x <= 491;
				I83x <= 753;
				I84x <= 1403;
				I85x <= 547;
				I86x <= 0;
				I87x <= 0;
				I88x <= 0;
				I89x <= 0;
				I90x <= 0;
				I91x <= 0;
				I92x <= 0;
				I93x <= 0;
				I94x <= 0;
				I95x <= 0;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01100000:begin
				I0x <= 8192;
				I1x <= 5427;
				I2x <= 4265;
				I3x <= 3611;
				I4x <= 2809;
				I5x <= 1173;
				I6x <= 1712;
				I7x <= 2687;
				I8x <= 2302;
				I9x <= 1238;
				I10x <= 1231;
				I11x <= 1353;
				I12x <= 1372;
				I13x <= 1481;
				I14x <= 1475;
				I15x <= 1539;
				I16x <= 1507;
				I17x <= 1539;
				I18x <= 1565;
				I19x <= 1578;
				I20x <= 1571;
				I21x <= 1648;
				I22x <= 1642;
				I23x <= 1699;
				I24x <= 1635;
				I25x <= 1629;
				I26x <= 1693;
				I27x <= 1770;
				I28x <= 1809;
				I29x <= 1892;
				I30x <= 1937;
				I31x <= 1924;
				I32x <= 1886;
				I33x <= 1879;
				I34x <= 1873;
				I35x <= 1809;
				I36x <= 1764;
				I37x <= 1655;
				I38x <= 1513;
				I39x <= 1411;
				I40x <= 1334;
				I41x <= 1359;
				I42x <= 1488;
				I43x <= 1340;
				I44x <= 1347;
				I45x <= 1321;
				I46x <= 1372;
				I47x <= 1372;
				I48x <= 1340;
				I49x <= 1462;
				I50x <= 1424;
				I51x <= 1526;
				I52x <= 1699;
				I53x <= 1655;
				I54x <= 1642;
				I55x <= 1687;
				I56x <= 1661;
				I57x <= 1597;
				I58x <= 1635;
				I59x <= 1674;
				I60x <= 1616;
				I61x <= 1623;
				I62x <= 1488;
				I63x <= 1629;
				I64x <= 1597;
				I65x <= 1623;
				I66x <= 1488;
				I67x <= 1571;
				I68x <= 1597;
				I69x <= 1501;
				I70x <= 1398;
				I71x <= 1321;
				I72x <= 1250;
				I73x <= 1417;
				I74x <= 1385;
				I75x <= 1424;
				I76x <= 1379;
				I77x <= 1385;
				I78x <= 1321;
				I79x <= 1359;
				I80x <= 1308;
				I81x <= 1424;
				I82x <= 1552;
				I83x <= 1353;
				I84x <= 1398;
				I85x <= 1417;
				I86x <= 1353;
				I87x <= 1347;
				I88x <= 1353;
				I89x <= 1436;
				I90x <= 1462;
				I91x <= 1263;
				I92x <= 1308;
				I93x <= 1327;
				I94x <= 1392;
				I95x <= 1430;
				I96x <= 1443;
				I97x <= 1334;
				I98x <= 1353;
				I99x <= 1372;
				I100x <= 1424;
				I101x <= 1417;
				I102x <= 1469;
				I103x <= 1443;
				I104x <= 1379;
				I105x <= 1302;
				I106x <= 1443;
				I107x <= 1539;
				I108x <= 2155;
				I109x <= 2527;
				I110x <= 2796;
				I111x <= 3092;
				I112x <= 3630;
				I113x <= 4272;
				I114x <= 4650;
				I115x <= 4792;
				I116x <= 4529;
				I117x <= 3451;
				I118x <= 2072;
				I119x <= 1738;
				I120x <= 1526;
				I121x <= 1494;
				I122x <= 1430;
				I123x <= 1424;
				I124x <= 1327;
				I125x <= 1289;
				I126x <= 1244;
				I127x <= 102;
				I128x <= 0;
				I129x <= 1911;
				I130x <= 6652;
				I131x <= 7736;
				I132x <= 5067;
				I133x <= 4265;
				I134x <= 3714;
				I135x <= 2149;
				I136x <= 1167;
				I137x <= 2559;
				I138x <= 2752;
				I139x <= 2123;
				I140x <= 1616;
				I141x <= 1648;
				I142x <= 1648;
				I143x <= 1706;
				I144x <= 1642;
				I145x <= 1783;
				I146x <= 1815;
				I147x <= 1969;
				I148x <= 1860;
				I149x <= 1886;
				I150x <= 1924;
				I151x <= 1898;
				I152x <= 1969;
				I153x <= 2181;
				I154x <= 2174;
				I155x <= 2136;
				I156x <= 2174;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01100001:begin
				I0x <= 8128;
				I1x <= 6098;
				I2x <= 3079;
				I3x <= 1347;
				I4x <= 775;
				I5x <= 711;
				I6x <= 779;
				I7x <= 613;
				I8x <= 481;
				I9x <= 463;
				I10x <= 730;
				I11x <= 662;
				I12x <= 587;
				I13x <= 632;
				I14x <= 722;
				I15x <= 734;
				I16x <= 606;
				I17x <= 775;
				I18x <= 790;
				I19x <= 696;
				I20x <= 892;
				I21x <= 1008;
				I22x <= 971;
				I23x <= 1065;
				I24x <= 1140;
				I25x <= 1216;
				I26x <= 1366;
				I27x <= 1584;
				I28x <= 1528;
				I29x <= 1600;
				I30x <= 1878;
				I31x <= 1863;
				I32x <= 1871;
				I33x <= 1927;
				I34x <= 1867;
				I35x <= 1859;
				I36x <= 1848;
				I37x <= 1626;
				I38x <= 1344;
				I39x <= 1174;
				I40x <= 1170;
				I41x <= 914;
				I42x <= 700;
				I43x <= 843;
				I44x <= 662;
				I45x <= 628;
				I46x <= 775;
				I47x <= 816;
				I48x <= 606;
				I49x <= 700;
				I50x <= 737;
				I51x <= 715;
				I52x <= 711;
				I53x <= 719;
				I54x <= 707;
				I55x <= 719;
				I56x <= 734;
				I57x <= 719;
				I58x <= 640;
				I59x <= 700;
				I60x <= 715;
				I61x <= 606;
				I62x <= 692;
				I63x <= 666;
				I64x <= 515;
				I65x <= 564;
				I66x <= 704;
				I67x <= 715;
				I68x <= 500;
				I69x <= 598;
				I70x <= 572;
				I71x <= 542;
				I72x <= 692;
				I73x <= 628;
				I74x <= 564;
				I75x <= 730;
				I76x <= 824;
				I77x <= 990;
				I78x <= 907;
				I79x <= 1189;
				I80x <= 1264;
				I81x <= 1362;
				I82x <= 1532;
				I83x <= 1581;
				I84x <= 1295;
				I85x <= 1167;
				I86x <= 896;
				I87x <= 621;
				I88x <= 417;
				I89x <= 335;
				I90x <= 402;
				I91x <= 361;
				I92x <= 455;
				I93x <= 353;
				I94x <= 244;
				I95x <= 308;
				I96x <= 380;
				I97x <= 308;
				I98x <= 0;
				I99x <= 380;
				I100x <= 1351;
				I101x <= 4487;
				I102x <= 8192;
				I103x <= 5963;
				I104x <= 2872;
				I105x <= 1189;
				I106x <= 771;
				I107x <= 609;
				I108x <= 391;
				I109x <= 429;
				I110x <= 395;
				I111x <= 376;
				I112x <= 425;
				I113x <= 335;
				I114x <= 240;
				I115x <= 519;
				I116x <= 466;
				I117x <= 500;
				I118x <= 523;
				I119x <= 493;
				I120x <= 628;
				I121x <= 677;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01100010:begin
				I0x <= 8192;
				I1x <= 4973;
				I2x <= 3703;
				I3x <= 1447;
				I4x <= 974;
				I5x <= 931;
				I6x <= 1065;
				I7x <= 979;
				I8x <= 1060;
				I9x <= 1092;
				I10x <= 1119;
				I11x <= 1108;
				I12x <= 1211;
				I13x <= 1237;
				I14x <= 1221;
				I15x <= 1259;
				I16x <= 1415;
				I17x <= 1415;
				I18x <= 1501;
				I19x <= 1539;
				I20x <= 1609;
				I21x <= 1647;
				I22x <= 1733;
				I23x <= 1883;
				I24x <= 1932;
				I25x <= 2013;
				I26x <= 2126;
				I27x <= 2163;
				I28x <= 2314;
				I29x <= 2282;
				I30x <= 2196;
				I31x <= 2109;
				I32x <= 1948;
				I33x <= 1754;
				I34x <= 1598;
				I35x <= 1431;
				I36x <= 1345;
				I37x <= 1324;
				I38x <= 1383;
				I39x <= 1394;
				I40x <= 1356;
				I41x <= 1350;
				I42x <= 1372;
				I43x <= 1377;
				I44x <= 1388;
				I45x <= 1442;
				I46x <= 1507;
				I47x <= 1582;
				I48x <= 1501;
				I49x <= 1555;
				I50x <= 1501;
				I51x <= 1533;
				I52x <= 1469;
				I53x <= 1523;
				I54x <= 1474;
				I55x <= 1377;
				I56x <= 1404;
				I57x <= 1442;
				I58x <= 1426;
				I59x <= 1464;
				I60x <= 1722;
				I61x <= 2072;
				I62x <= 2190;
				I63x <= 2287;
				I64x <= 2271;
				I65x <= 2255;
				I66x <= 1835;
				I67x <= 1813;
				I68x <= 1399;
				I69x <= 1162;
				I70x <= 1194;
				I71x <= 1054;
				I72x <= 1017;
				I73x <= 1060;
				I74x <= 1065;
				I75x <= 974;
				I76x <= 457;
				I77x <= 0;
				I78x <= 2325;
				I79x <= 7266;
				I80x <= 7944;
				I81x <= 3805;
				I82x <= 2029;
				I83x <= 1291;
				I84x <= 1162;
				I85x <= 1394;
				I86x <= 1329;
				I87x <= 1297;
				I88x <= 1350;
				I89x <= 1291;
				I90x <= 1340;
				I91x <= 1431;
				I92x <= 1544;
				I93x <= 1544;
				I94x <= 1533;
				I95x <= 1571;
				I96x <= 0;
				I97x <= 0;
				I98x <= 0;
				I99x <= 0;
				I100x <= 0;
				I101x <= 0;
				I102x <= 0;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

			9b'0b01100011:begin
				I0x <= 8192;
				I1x <= 7478;
				I2x <= 7260;
				I3x <= 7147;
				I4x <= 7249;
				I5x <= 5519;
				I6x <= 3853;
				I7x <= 2584;
				I8x <= 1824;
				I9x <= 1687;
				I10x <= 1374;
				I11x <= 1262;
				I12x <= 1321;
				I13x <= 1198;
				I14x <= 1132;
				I15x <= 1111;
				I16x <= 1068;
				I17x <= 907;
				I18x <= 798;
				I19x <= 769;
				I20x <= 791;
				I21x <= 755;
				I22x <= 534;
				I23x <= 527;
				I24x <= 326;
				I25x <= 151;
				I26x <= 414;
				I27x <= 144;
				I28x <= 203;
				I29x <= 49;
				I30x <= 0;
				I31x <= 418;
				I32x <= 326;
				I33x <= 541;
				I34x <= 513;
				I35x <= 938;
				I36x <= 1357;
				I37x <= 1508;
				I38x <= 1909;
				I39x <= 1968;
				I40x <= 2320;
				I41x <= 2362;
				I42x <= 2106;
				I43x <= 2309;
				I44x <= 2039;
				I45x <= 2267;
				I46x <= 2218;
				I47x <= 2070;
				I48x <= 2063;
				I49x <= 1884;
				I50x <= 2039;
				I51x <= 2067;
				I52x <= 1831;
				I53x <= 2042;
				I54x <= 1944;
				I55x <= 1940;
				I56x <= 1842;
				I57x <= 1641;
				I58x <= 1659;
				I59x <= 1779;
				I60x <= 1729;
				I61x <= 1993;
				I62x <= 2338;
				I63x <= 2738;
				I64x <= 3157;
				I65x <= 3480;
				I66x <= 3793;
				I67x <= 3828;
				I68x <= 3804;
				I69x <= 3635;
				I70x <= 3069;
				I71x <= 2974;
				I72x <= 2334;
				I73x <= 2158;
				I74x <= 1965;
				I75x <= 1687;
				I76x <= 2000;
				I77x <= 2144;
				I78x <= 2598;
				I79x <= 3656;
				I80x <= 4060;
				I81x <= 4292;
				I82x <= 4584;
				I83x <= 6149;
				I84x <= 5716;
				I85x <= 6332;
				I86x <= 5720;
				I87x <= 5948;
				I88x <= 6321;
				I89x <= 6117;
				I90x <= 4595;
				I91x <= 3167;
				I92x <= 1975;
				I93x <= 1241;
				I94x <= 1223;
				I95x <= 1139;
				I96x <= 1153;
				I97x <= 956;
				I98x <= 1075;
				I99x <= 1128;
				I100x <= 1058;
				I101x <= 1047;
				I102x <= 857;
				I103x <= 0;
				I104x <= 0;
				I105x <= 0;
				I106x <= 0;
				I107x <= 0;
				I108x <= 0;
				I109x <= 0;
				I110x <= 0;
				I111x <= 0;
				I112x <= 0;
				I113x <= 0;
				I114x <= 0;
				I115x <= 0;
				I116x <= 0;
				I117x <= 0;
				I118x <= 0;
				I119x <= 0;
				I120x <= 0;
				I121x <= 0;
				I122x <= 0;
				I123x <= 0;
				I124x <= 0;
				I125x <= 0;
				I126x <= 0;
				I127x <= 0;
				I128x <= 0;
				I129x <= 0;
				I130x <= 0;
				I131x <= 0;
				I132x <= 0;
				I133x <= 0;
				I134x <= 0;
				I135x <= 0;
				I136x <= 0;
				I137x <= 0;
				I138x <= 0;
				I139x <= 0;
				I140x <= 0;
				I141x <= 0;
				I142x <= 0;
				I143x <= 0;
				I144x <= 0;
				I145x <= 0;
				I146x <= 0;
				I147x <= 0;
				I148x <= 0;
				I149x <= 0;
				I150x <= 0;
				I151x <= 0;
				I152x <= 0;
				I153x <= 0;
				I154x <= 0;
				I155x <= 0;
				I156x <= 0;
				I157x <= 0;
				I158x <= 0;
				I159x <= 0;
				I160x <= 0;
				I161x <= 0;
				I162x <= 0;
				I163x <= 0;
				I164x <= 0;
				I165x <= 0;
				I166x <= 0;
				I167x <= 0;
				I168x <= 0;
				I169x <= 0;
				I170x <= 0;
				I171x <= 0;
				I172x <= 0;
				I173x <= 0;
				I174x <= 0;
				I175x <= 0;
				I176x <= 0;
				I177x <= 0;
				I178x <= 0;
				I179x <= 0;
				I180x <= 0;
				I181x <= 0;
				I182x <= 0;
				I183x <= 0;
				I184x <= 0;
				I185x <= 0;
				I186x <= 0;
			end

		endcase
	end
endmodule
