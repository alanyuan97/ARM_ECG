module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = -1052;
	I1x = 8041;
	I2x = 1403;
	I3x = 7197;
	I4x = 3283;
	I5x = 6732;
	I6x = -6935;
	I7x = -1872;
	I8x = 7366;
	I9x = -362;
	I10x = 2189;
	I11x = 3216;
	I12x = 3623;
	I13x = 7155;
	I14x = 935;
	I15x = 543;
	I16x = 7990;
	I17x = 5797;
	I18x = 6436;
	I19x = 631;
	I20x = -640;
	I21x = 5604;
	I22x = -3323;
	I23x = -5846;
	I24x = -4997;
	I25x = 1368;
	I26x = 1359;
	I27x = 2788;
	I28x = -4161;
	I29x = 3396;
	I30x = -3533;
	I31x = -4398;
	I32x = 7818;
	I33x = -5696;
	I34x = -3661;
	I35x = 2611;
	I36x = -1270;
	I37x = 6727;
	I38x = -2390;
	I39x = 6079;
	I40x = -1436;
	I41x = 4564;
	I42x = 1508;
	I43x = 511;
	I44x = 3479;
	I45x = -169;
	I46x = 5522;
	I47x = -981;
	I48x = -6558;
	I49x = -11;
	I50x = 4978;
	I51x = -704;
	I52x = -409;
	I53x = -6474;
	I54x = 3623;
	I55x = 7759;
	I56x = -6735;
	I57x = -6485;
	I58x = -4745;
	I59x = 3256;
	I60x = 1922;
	I61x = -4971;
	I62x = -4366;
	I63x = -2349;
	I64x = -7212;
	I65x = -2747;
	I66x = -3049;
	I67x = -2004;
	I68x = 7756;
	I69x = 1040;
	I70x = 3309;
	I71x = -7814;
	I72x = -6714;
	I73x = -1647;
	I74x = 1919;
	I75x = -1006;
	I76x = -6332;
	I77x = -953;
	I78x = -5241;
	I79x = -159;
	I80x = 4606;
	I81x = 7138;
	I82x = -6424;
	I83x = -6914;
	I84x = 4852;
	I85x = -1427;
	I86x = 6750;
	I87x = 166;
	I88x = -2937;
	I89x = 372;
	I90x = -4661;
	I91x = 5264;
	I92x = 5843;
	I93x = -1891;
	I94x = -5072;
	I95x = 2652;
	I96x = -5906;
	I97x = -1334;
	I98x = -1643;
	I99x = 3039;
	I100x = -326;
	I101x = -5403;
	I102x = 5611;
	I103x = 3012;
	I104x = 8123;
	I105x = -1291;
	I106x = -4691;
	I107x = -6469;
	I108x = 7246;
	I109x = 1918;
	I110x = -1560;
	I111x = 5314;
	I112x = -258;
	I113x = -999;
	I114x = -7230;
	I115x = -698;
	I116x = -6918;
	I117x = -4042;
	I118x = -7706;
	I119x = 8037;
	I120x = 3951;
	I121x = -621;
	I122x = 6238;
	I123x = 325;
	I124x = 6052;
	I125x = -8158;
	I126x = 6614;
	I127x = -6883;
	I128x = 6932;
	I129x = 4143;
	I130x = 5286;
	I131x = 1087;
	I132x = 4437;
	I133x = -7503;
	I134x = 8105;
	I135x = 6127;
	I136x = -1033;
	I137x = 5787;
	I138x = -6044;
	I139x = -2644;
	I140x = -7643;
	I141x = -1385;
	I142x = 608;
	I143x = 5940;
	I144x = 469;
	I145x = 5386;
	I146x = 6927;
	I147x = 7112;
	I148x = -437;
	I149x = 7991;
	I150x = -5105;
	I151x = -995;
	I152x = -2001;
	I153x = 1784;
	I154x = 5403;
	I155x = -4923;
	I156x = 1526;
	I157x = -215;
	I158x = -7105;
	I159x = -2787;
	I160x = 8053;
	I161x = 2323;
	I162x = -4894;
	I163x = 1823;
	I164x = 4281;
	I165x = -2601;
	I166x = -5247;
	I167x = 4171;
	I168x = -2071;
	I169x = 1819;
	I170x = 5697;
	I171x = -2894;
	I172x = -2227;
	I173x = -2215;
	I174x = 1795;
	I175x = 6506;
	I176x = -461;
	I177x = 1274;
	I178x = 5910;
	I179x = 195;
	I180x = 3624;
	I181x = 2752;
	I182x = -1291;
	I183x = 4924;
	I184x = 632;
	I185x = -5298;
	I186x = 7394;
	end
endmodule
[0.         3.07167073 0.         0.         0.        ] 

 [0, 25163, 0, 0, 0] 

 ['0000000000000000', '0110001001001011', '0000000000000000', '0000000000000000', '0000000000000000']
