module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 41;
	I1x = -33;
	I2x = 1;
	I3x = 38;
	I4x = 23;
	I5x = 59;
	I6x = -40;
	I7x = 18;
	I8x = 9;
	I9x = -54;
	I10x = -9;
	I11x = 25;
	I12x = 37;
	I13x = 37;
	I14x = -17;
	I15x = 12;
	I16x = 34;
	I17x = -36;
	I18x = -25;
	I19x = -13;
	I20x = 56;
	I21x = -24;
	I22x = 17;
	I23x = -50;
	I24x = 3;
	I25x = 24;
	I26x = -59;
	I27x = 62;
	I28x = 46;
	I29x = -10;
	I30x = 46;
	I31x = -43;
	I32x = -61;
	I33x = 12;
	I34x = 5;
	I35x = -24;
	I36x = 26;
	I37x = -44;
	I38x = 40;
	I39x = -12;
	I40x = 60;
	I41x = 6;
	I42x = 4;
	I43x = 61;
	I44x = 41;
	I45x = -63;
	I46x = -14;
	I47x = 36;
	I48x = -22;
	I49x = 27;
	I50x = -34;
	I51x = -11;
	I52x = -17;
	I53x = -6;
	I54x = -52;
	I55x = -26;
	I56x = 49;
	I57x = 40;
	I58x = -23;
	I59x = -48;
	I60x = 14;
	I61x = 32;
	I62x = -40;
	I63x = -7;
	I64x = -27;
	I65x = 20;
	I66x = 42;
	I67x = -12;
	I68x = 28;
	I69x = 28;
	I70x = -47;
	I71x = 52;
	I72x = 9;
	I73x = 60;
	I74x = -62;
	I75x = 8;
	I76x = -46;
	I77x = 34;
	I78x = -53;
	I79x = -60;
	I80x = -24;
	I81x = 60;
	I82x = -57;
	I83x = -40;
	I84x = -28;
	I85x = 35;
	I86x = 21;
	I87x = 61;
	I88x = -30;
	I89x = 1;
	I90x = -43;
	I91x = -53;
	I92x = 2;
	I93x = 9;
	I94x = 26;
	I95x = -34;
	I96x = -4;
	I97x = 28;
	I98x = 29;
	I99x = 50;
	I100x = 50;
	I101x = -37;
	I102x = -20;
	I103x = 61;
	I104x = -5;
	I105x = 15;
	I106x = -55;
	I107x = 14;
	I108x = 32;
	I109x = -25;
	I110x = -53;
	I111x = -6;
	I112x = 17;
	I113x = -39;
	I114x = -48;
	I115x = 41;
	I116x = -42;
	I117x = -38;
	I118x = 39;
	I119x = -59;
	I120x = -45;
	I121x = 0;
	I122x = 25;
	I123x = 10;
	I124x = 26;
	I125x = -2;
	I126x = 5;
	I127x = 7;
	I128x = -29;
	I129x = -22;
	I130x = -10;
	I131x = 58;
	I132x = -61;
	I133x = 60;
	I134x = -15;
	I135x = -22;
	I136x = -39;
	I137x = 61;
	I138x = 12;
	I139x = 22;
	I140x = 18;
	I141x = 8;
	I142x = -39;
	I143x = -50;
	I144x = 17;
	I145x = 11;
	I146x = -3;
	I147x = 35;
	I148x = 34;
	I149x = 53;
	I150x = -63;
	I151x = 28;
	I152x = -1;
	I153x = 0;
	I154x = -43;
	I155x = 11;
	I156x = 47;
	I157x = -56;
	I158x = -25;
	I159x = -45;
	I160x = -45;
	I161x = 52;
	I162x = 45;
	I163x = 56;
	I164x = 27;
	I165x = -48;
	I166x = -13;
	I167x = -11;
	I168x = 13;
	I169x = 61;
	I170x = 5;
	I171x = 0;
	I172x = 32;
	I173x = -4;
	I174x = 35;
	I175x = -5;
	I176x = -23;
	I177x = 54;
	I178x = -28;
	I179x = 58;
	I180x = 14;
	I181x = 47;
	I182x = 45;
	I183x = 57;
	I184x = -14;
	I185x = -1;
	I186x = -4;
	end
endmodule
 

