module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	output [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	input EN;
	
	always@(EN)
	begin
	I0x = 32'b00111111011111110111110011101110;
	I1x = 32'b00111111000100111011011001000110;
	I2x = 32'b00111110101101011100001010001111;
	I3x = 32'b00111110001001011110001101010100;
	I4x = 32'b00111110001000111101011100001010;
	I5x = 32'b00111110001100110011001100110011;
	I6x = 32'b00111110001101010011111101111101;
	I7x = 32'b00111110001011010000111001010110;
	I8x = 32'b00111110001100100010110100001110;
	I9x = 32'b00111110001011010000111001010110;
	I10x = 32'b00111110001010110000001000001100;
	I11x = 32'b00111110001011110001101010100000;
	I12x = 32'b00111110001011110001101010100000;
	I13x = 32'b00111110001101010011111101111101;
	I14x = 32'b00111110001100100010110100001110;
	I15x = 32'b00111110001100110011001100110011;
	I16x = 32'b00111110001111000110101001111111;
	I17x = 32'b00111110010000001000001100010010;
	I18x = 32'b00111110010011001100110011001101;
	I19x = 32'b00111110010011111101111100111011;
	I20x = 32'b00111110010101100000010000011001;
	I21x = 32'b00111110011001010110000001000010;
	I22x = 32'b00111110011011111001110110110010;
	I23x = 32'b00111110100000011000100100110111;
	I24x = 32'b00111110100001101010011111110000;
	I25x = 32'b00111110100011010100111111011111;
	I26x = 32'b00111110100101111000110101010000;
	I27x = 32'b00111110100111000010100011110110;
	I28x = 32'b00111110101001000101101000011101;
	I29x = 32'b00111110101001011110001101010100;
	I30x = 32'b00111110101010001111010111000011;
	I31x = 32'b00111110101011001000101101000100;
	I32x = 32'b00111110101001101110100101111001;
	I33x = 32'b00111110101000000100000110001001;
	I34x = 32'b00111110100011101101100100010111;
	I35x = 32'b00111110100000011000100100110111;
	I36x = 32'b00111110011011101001011110001101;
	I37x = 32'b00111110010101100000010000011001;
	I38x = 32'b00111110010011001100110011001101;
	I39x = 32'b00111110001111000110101001111111;
	I40x = 32'b00111110001101000011100101011000;
	I41x = 32'b00111110001101000011100101011000;
	I42x = 32'b00111110001100000010000011000101;
	I43x = 32'b00111110001101000011100101011000;
	I44x = 32'b00111110001011100001010001111011;
	I45x = 32'b00111110001011000000100000110001;
	I46x = 32'b00111110001011110001101010100000;
	I47x = 32'b00111110001011010000111001010110;
	I48x = 32'b00111110001101010011111101111101;
	I49x = 32'b00111110001100000010000011000101;
	I50x = 32'b00111110001011110001101010100000;
	I51x = 32'b00111110001100000010000011000101;
	I52x = 32'b00111110001011110001101010100000;
	I53x = 32'b00111110001101100100010110100010;
	I54x = 32'b00111110001100000010000011000101;
	I55x = 32'b00111110001011110001101010100000;
	I56x = 32'b00111110001100100010110100001110;
	I57x = 32'b00111110001011110001101010100000;
	I58x = 32'b00111110001101010011111101111101;
	I59x = 32'b00111110001011100001010001111011;
	I60x = 32'b00111110001010011111101111100111;
	I61x = 32'b00111110001010011111101111100111;
	I62x = 32'b00111110001001111110111110011110;
	I63x = 32'b00111110001011000000100000110001;
	I64x = 32'b00111110001001001101110100101111;
	I65x = 32'b00111110001000101101000011100101;
	I66x = 32'b00111110001001011110001101010100;
	I67x = 32'b00111110001000111101011100001010;
	I68x = 32'b00111110001010011111101111100111;
	I69x = 32'b00111110001001001101110100101111;
	I70x = 32'b00111110001001101110100101111001;
	I71x = 32'b00111110001110010101100000010000;
	I72x = 32'b00111110010000011000100100110111;
	I73x = 32'b00111110010011101101100100010111;
	I74x = 32'b00111110010001011010000111001011;
	I75x = 32'b00111110010010011011101001011110;
	I76x = 32'b00111110010101110000101000111101;
	I77x = 32'b00111110010111000010100011110110;
	I78x = 32'b00111110010111110011101101100100;
	I79x = 32'b00111110010011011101001011110010;
	I80x = 32'b00111110001100000010000011000101;
	I81x = 32'b00111110001000111101011100001010;
	I82x = 32'b00111110000110101001111110111110;
	I83x = 32'b00111110000110101001111110111110;
	I84x = 32'b00111110000011110101110000101001;
	I85x = 32'b00111110000010100011110101110001;
	I86x = 32'b00111110000011010100111111011111;
	I87x = 32'b00111110000010000011000100100111;
	I88x = 32'b00111110000011110101110000101001;
	I89x = 32'b00111110000010110100001110010110;
	I90x = 32'b00111110000010010011011101001100;
	I91x = 32'b00111110000010100011110101110001;
	I92x = 32'b00111101111011111001110110110010;
	I93x = 32'b00000000000000000000000000000000;
	I94x = 32'b00111100101001010111101001111000;
	I95x = 32'b00111110011101101100100010110100;
	I96x = 32'b00111111000111001110110110010001;
	I97x = 32'b00111111100000000000000000000000;
	I98x = 32'b00111111001011010100111111011111;
	I99x = 32'b00111110110110000001000001100010;
	I100x = 32'b00111110010011001100110011001101;
	I101x = 32'b00111110000101101000011100101011;
	I102x = 32'b00111110001011010000111001010110;
	I103x = 32'b00111110001110000101000111101100;
	I104x = 32'b00111110001001001101110100101111;
	I105x = 32'b00111110001001001101110100101111;
	I106x = 32'b00111110001001111110111110011110;
	I107x = 32'b00111110001001101110100101111001;
	I108x = 32'b00111110001011110001101010100000;
	I109x = 32'b00111110001011010000111001010110;
	I110x = 32'b00111110001100010010011011101001;
	I111x = 32'b00111110001110010101100000010000;
	I112x = 32'b00111110001110010101100000010000;
	I113x = 32'b00111110010000011000100100110111;
	I114x = 32'b00111110010000011000100100110111;
	I115x = 32'b00000000000000000000000000000000;
	I116x = 32'b00000000000000000000000000000000;
	I117x = 32'b00000000000000000000000000000000;
	I118x = 32'b00000000000000000000000000000000;
	I119x = 32'b00000000000000000000000000000000;
	I120x = 32'b00000000000000000000000000000000;
	I121x = 32'b00000000000000000000000000000000;
	I122x = 32'b00000000000000000000000000000000;
	I123x = 32'b00000000000000000000000000000000;
	I124x = 32'b00000000000000000000000000000000;
	I125x = 32'b00000000000000000000000000000000;
	I126x = 32'b00000000000000000000000000000000;
	I127x = 32'b00000000000000000000000000000000;
	I128x = 32'b00000000000000000000000000000000;
	I129x = 32'b00000000000000000000000000000000;
	I130x = 32'b00000000000000000000000000000000;
	I131x = 32'b00000000000000000000000000000000;
	I132x = 32'b00000000000000000000000000000000;
	I133x = 32'b00000000000000000000000000000000;
	I134x = 32'b00000000000000000000000000000000;
	I135x = 32'b00000000000000000000000000000000;
	I136x = 32'b00000000000000000000000000000000;
	I137x = 32'b00000000000000000000000000000000;
	I138x = 32'b00000000000000000000000000000000;
	I139x = 32'b00000000000000000000000000000000;
	I140x = 32'b00000000000000000000000000000000;
	I141x = 32'b00000000000000000000000000000000;
	I142x = 32'b00000000000000000000000000000000;
	I143x = 32'b00000000000000000000000000000000;
	I144x = 32'b00000000000000000000000000000000;
	I145x = 32'b00000000000000000000000000000000;
	I146x = 32'b00000000000000000000000000000000;
	I147x = 32'b00000000000000000000000000000000;
	I148x = 32'b00000000000000000000000000000000;
	I149x = 32'b00000000000000000000000000000000;
	I150x = 32'b00000000000000000000000000000000;
	I151x = 32'b00000000000000000000000000000000;
	I152x = 32'b00000000000000000000000000000000;
	I153x = 32'b00000000000000000000000000000000;
	I154x = 32'b00000000000000000000000000000000;
	I155x = 32'b00000000000000000000000000000000;
	I156x = 32'b00000000000000000000000000000000;
	I157x = 32'b00000000000000000000000000000000;
	I158x = 32'b00000000000000000000000000000000;
	I159x = 32'b00000000000000000000000000000000;
	I160x = 32'b00000000000000000000000000000000;
	I161x = 32'b00000000000000000000000000000000;
	I162x = 32'b00000000000000000000000000000000;
	I163x = 32'b00000000000000000000000000000000;
	I164x = 32'b00000000000000000000000000000000;
	I165x = 32'b00000000000000000000000000000000;
	I166x = 32'b00000000000000000000000000000000;
	I167x = 32'b00000000000000000000000000000000;
	I168x = 32'b00000000000000000000000000000000;
	I169x = 32'b00000000000000000000000000000000;
	I170x = 32'b00000000000000000000000000000000;
	I171x = 32'b00000000000000000000000000000000;
	I172x = 32'b00000000000000000000000000000000;
	I173x = 32'b00000000000000000000000000000000;
	I174x = 32'b00000000000000000000000000000000;
	I175x = 32'b00000000000000000000000000000000;
	I176x = 32'b00000000000000000000000000000000;
	I177x = 32'b00000000000000000000000000000000;
	I178x = 32'b00000000000000000000000000000000;
	I179x = 32'b00000000000000000000000000000000;
	I180x = 32'b00000000000000000000000000000000;
	I181x = 32'b00000000000000000000000000000000;
	I182x = 32'b00000000000000000000000000000000;
	I183x = 32'b00000000000000000000000000000000;
	I184x = 32'b00000000000000000000000000000000;
	I185x = 32'b00000000000000000000000000000000;
	I186x = 32'b00000000000000000000000000000000;
	end
endmodule
