module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 8192;
	I1x = 6579;
	I2x = 1825;
	I3x = 160;
	I4x = 808;
	I5x = 1090;
	I6x = 851;
	I7x = 1043;
	I8x = 1160;
	I9x = 1029;
	I10x = 1412;
	I11x = 1277;
	I12x = 1390;
	I13x = 1373;
	I14x = 1221;
	I15x = 1525;
	I16x = 1403;
	I17x = 1516;
	I18x = 1503;
	I19x = 1368;
	I20x = 1664;
	I21x = 1529;
	I22x = 1612;
	I23x = 1655;
	I24x = 1503;
	I25x = 1868;
	I26x = 1833;
	I27x = 1929;
	I28x = 1968;
	I29x = 1816;
	I30x = 2203;
	I31x = 2081;
	I32x = 2094;
	I33x = 2059;
	I34x = 1877;
	I35x = 2146;
	I36x = 1929;
	I37x = 1899;
	I38x = 1799;
	I39x = 1538;
	I40x = 1816;
	I41x = 1720;
	I42x = 1716;
	I43x = 1703;
	I44x = 1442;
	I45x = 1781;
	I46x = 1664;
	I47x = 1655;
	I48x = 1590;
	I49x = 1386;
	I50x = 1681;
	I51x = 1555;
	I52x = 1534;
	I53x = 1581;
	I54x = 1360;
	I55x = 1690;
	I56x = 1547;
	I57x = 1629;
	I58x = 1642;
	I59x = 1438;
	I60x = 1699;
	I61x = 1612;
	I62x = 1581;
	I63x = 1603;
	I64x = 1381;
	I65x = 1660;
	I66x = 1547;
	I67x = 1547;
	I68x = 1647;
	I69x = 1464;
	I70x = 1825;
	I71x = 1755;
	I72x = 1864;
	I73x = 1946;
	I74x = 1773;
	I75x = 1973;
	I76x = 1942;
	I77x = 1838;
	I78x = 1664;
	I79x = 1029;
	I80x = 1477;
	I81x = 1403;
	I82x = 1529;
	I83x = 1547;
	I84x = 1190;
	I85x = 1421;
	I86x = 1573;
	I87x = 2520;
	I88x = 3972;
	I89x = 4558;
	I90x = 6675;
	I91x = 8131;
	I92x = 4915;
	I93x = 1038;
	I94x = 0;
	I95x = 1021;
	I96x = 756;
	I97x = 817;
	I98x = 969;
	I99x = 860;
	I100x = 1134;
	I101x = 1082;
	I102x = 1177;
	I103x = 1260;
	I104x = 1029;
	I105x = 1247;
	I106x = 1208;
	I107x = 1242;
	I108x = 1408;
	I109x = 0;
	I110x = 0;
	I111x = 0;
	I112x = 0;
	I113x = 0;
	I114x = 0;
	I115x = 0;
	I116x = 0;
	I117x = 0;
	I118x = 0;
	I119x = 0;
	I120x = 0;
	I121x = 0;
	I122x = 0;
	I123x = 0;
	I124x = 0;
	I125x = 0;
	I126x = 0;
	I127x = 0;
	I128x = 0;
	I129x = 0;
	I130x = 0;
	I131x = 0;
	I132x = 0;
	I133x = 0;
	I134x = 0;
	I135x = 0;
	I136x = 0;
	I137x = 0;
	I138x = 0;
	I139x = 0;
	I140x = 0;
	I141x = 0;
	I142x = 0;
	I143x = 0;
	I144x = 0;
	I145x = 0;
	I146x = 0;
	I147x = 0;
	I148x = 0;
	I149x = 0;
	I150x = 0;
	I151x = 0;
	I152x = 0;
	I153x = 0;
	I154x = 0;
	I155x = 0;
	I156x = 0;
	I157x = 0;
	I158x = 0;
	I159x = 0;
	I160x = 0;
	I161x = 0;
	I162x = 0;
	I163x = 0;
	I164x = 0;
	I165x = 0;
	I166x = 0;
	I167x = 0;
	I168x = 0;
	I169x = 0;
	I170x = 0;
	I171x = 0;
	I172x = 0;
	I173x = 0;
	I174x = 0;
	I175x = 0;
	I176x = 0;
	I177x = 0;
	I178x = 0;
	I179x = 0;
	I180x = 0;
	I181x = 0;
	I182x = 0;
	I183x = 0;
	I184x = 0;
	I185x = 0;
	I186x = 0;
	end
endmodule
