module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = -6254;
	I1x = -6278;
	I2x = 1838;
	I3x = 3460;
	I4x = 6751;
	I5x = 6204;
	I6x = 5942;
	I7x = -7333;
	I8x = 6188;
	I9x = -6423;
	I10x = 5297;
	I11x = 5728;
	I12x = 4304;
	I13x = -3680;
	I14x = 5501;
	I15x = -4096;
	I16x = -799;
	I17x = 6798;
	I18x = -445;
	I19x = -6285;
	I20x = -6571;
	I21x = -7490;
	I22x = -6964;
	I23x = -3351;
	I24x = -3132;
	I25x = 6120;
	I26x = -6768;
	I27x = 3210;
	I28x = -1437;
	I29x = -1453;
	I30x = 3756;
	I31x = -3718;
	I32x = 7353;
	I33x = 5634;
	I34x = 3909;
	I35x = 6913;
	I36x = 3594;
	I37x = -7280;
	I38x = 5794;
	I39x = -4671;
	I40x = 1;
	I41x = 6207;
	I42x = 2844;
	I43x = -7711;
	I44x = -4057;
	I45x = -6984;
	I46x = 2922;
	I47x = -7380;
	I48x = -8187;
	I49x = 6977;
	I50x = 6873;
	I51x = 2803;
	I52x = 7592;
	I53x = 2091;
	I54x = 2381;
	I55x = -2761;
	I56x = 4074;
	I57x = -5907;
	I58x = -1583;
	I59x = 6123;
	I60x = 4894;
	I61x = -6041;
	I62x = -2769;
	I63x = -2485;
	I64x = -6700;
	I65x = -3925;
	I66x = 8184;
	I67x = 1172;
	I68x = 5572;
	I69x = -4460;
	I70x = -404;
	I71x = -3565;
	I72x = 5045;
	I73x = -5612;
	I74x = 508;
	I75x = -1804;
	I76x = 2288;
	I77x = -5333;
	I78x = -4151;
	I79x = 1813;
	I80x = -310;
	I81x = -3682;
	I82x = 6503;
	I83x = 6721;
	I84x = 4433;
	I85x = -3387;
	I86x = -1727;
	I87x = 4122;
	I88x = -7876;
	I89x = -2749;
	I90x = -2716;
	I91x = 3845;
	I92x = -7509;
	I93x = -5043;
	I94x = 1271;
	I95x = 1778;
	I96x = -5095;
	I97x = -145;
	I98x = -1537;
	I99x = 7004;
	I100x = 5918;
	I101x = 550;
	I102x = -5697;
	I103x = -7609;
	I104x = -7274;
	I105x = -7639;
	I106x = 8022;
	I107x = 6883;
	I108x = -2837;
	I109x = -5413;
	I110x = -2052;
	I111x = 4712;
	I112x = -2969;
	I113x = -5688;
	I114x = 3697;
	I115x = -7329;
	I116x = 6312;
	I117x = -7047;
	I118x = -772;
	I119x = -1977;
	I120x = 5123;
	I121x = 1057;
	I122x = 248;
	I123x = -630;
	I124x = -1120;
	I125x = -3766;
	I126x = -5471;
	I127x = -5661;
	I128x = 7827;
	I129x = 4636;
	I130x = 3244;
	I131x = 1996;
	I132x = 3274;
	I133x = 4695;
	I134x = 1962;
	I135x = -2558;
	I136x = 886;
	I137x = -5252;
	I138x = -4794;
	I139x = -7710;
	I140x = 4866;
	I141x = -2057;
	I142x = -7091;
	I143x = -5197;
	I144x = 4231;
	I145x = 3972;
	I146x = -409;
	I147x = -8010;
	I148x = -6800;
	I149x = -8150;
	I150x = -3294;
	I151x = 4471;
	I152x = 3824;
	I153x = -3212;
	I154x = -360;
	I155x = 519;
	I156x = 3261;
	I157x = -699;
	I158x = -6672;
	I159x = -7497;
	I160x = -724;
	I161x = -4085;
	I162x = 4539;
	I163x = 7405;
	I164x = 1146;
	I165x = 7955;
	I166x = -5902;
	I167x = -1414;
	I168x = -5498;
	I169x = -6079;
	I170x = 1348;
	I171x = 11;
	I172x = -2012;
	I173x = 6334;
	I174x = 7196;
	I175x = -1394;
	I176x = 2922;
	I177x = 6114;
	I178x = -891;
	I179x = 3858;
	I180x = 6204;
	I181x = 6035;
	I182x = -1437;
	I183x = -5701;
	I184x = 6978;
	I185x = -5560;
	I186x = -6306;
	end
endmodule
[0.         1.3739656  2.43033068 0.         0.71922951] 

 [0, 11255, 19909, 0, 5891] 

 ['0000000000000000', '0010101111110111', '0100110111000101', '0000000000000000', '0001011100000011']
