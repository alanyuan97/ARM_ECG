module rom_input(EN, clk, I0x, I1x, I2x, I3x, I4x, I5x, I6x, I7x, I8x, I9x, I10x, I11x, I12x, I13x, I14x, I15x, I16x, I17x, I18x, I19x, I20x, I21x, I22x, I23x, I24x, I25x, I26x, I27x, I28x, I29x, I30x, I31x, I32x, I33x, I34x, I35x, I36x, I37x, I38x, I39x, I40x, I41x, I42x, I43x, I44x, I45x, I46x, I47x, I48x, I49x, I50x, I51x, I52x, I53x, I54x, I55x, I56x, I57x, I58x, I59x, I60x, I61x, I62x, I63x, I64x, I65x, I66x, I67x, I68x, I69x, I70x, I71x, I72x, I73x, I74x, I75x, I76x, I77x, I78x, I79x, I80x, I81x, I82x, I83x, I84x, I85x, I86x, I87x, I88x, I89x, I90x, I91x, I92x, I93x, I94x, I95x, I96x, I97x, I98x, I99x, I100x, I101x, I102x, I103x, I104x, I105x, I106x, I107x, I108x, I109x, I110x, I111x, I112x, I113x, I114x, I115x, I116x, I117x, I118x, I119x, I120x, I121x, I122x, I123x, I124x, I125x, I126x, I127x, I128x, I129x, I130x, I131x, I132x, I133x, I134x, I135x, I136x, I137x, I138x, I139x, I140x, I141x, I142x, I143x, I144x, I145x, I146x, I147x, I148x, I149x, I150x, I151x, I152x, I153x, I154x, I155x, I156x, I157x, I158x, I159x, I160x, I161x, I162x, I163x, I164x, I165x, I166x, I167x, I168x, I169x, I170x, I171x, I172x, I173x, I174x, I175x, I176x, I177x, I178x, I179x, I180x, I181x, I182x, I183x, I184x, I185x, I186x);
	input EN, clk;
	output reg [7:0] I0x, I1x, I2x, I3x, I4x, I5x, I6x, I7x, I8x, I9x, I10x, I11x, I12x, I13x, I14x, I15x, I16x, I17x, I18x, I19x, I20x, I21x, I22x, I23x, I24x, I25x, I26x, I27x, I28x, I29x, I30x, I31x, I32x, I33x, I34x, I35x, I36x, I37x, I38x, I39x, I40x, I41x, I42x, I43x, I44x, I45x, I46x, I47x, I48x, I49x, I50x, I51x, I52x, I53x, I54x, I55x, I56x, I57x, I58x, I59x, I60x, I61x, I62x, I63x, I64x, I65x, I66x, I67x, I68x, I69x, I70x, I71x, I72x, I73x, I74x, I75x, I76x, I77x, I78x, I79x, I80x, I81x, I82x, I83x, I84x, I85x, I86x, I87x, I88x, I89x, I90x, I91x, I92x, I93x, I94x, I95x, I96x, I97x, I98x, I99x, I100x, I101x, I102x, I103x, I104x, I105x, I106x, I107x, I108x, I109x, I110x, I111x, I112x, I113x, I114x, I115x, I116x, I117x, I118x, I119x, I120x, I121x, I122x, I123x, I124x, I125x, I126x, I127x, I128x, I129x, I130x, I131x, I132x, I133x, I134x, I135x, I136x, I137x, I138x, I139x, I140x, I141x, I142x, I143x, I144x, I145x, I146x, I147x, I148x, I149x, I150x, I151x, I152x, I153x, I154x, I155x, I156x, I157x, I158x, I159x, I160x, I161x, I162x, I163x, I164x, I165x, I166x, I167x, I168x, I169x, I170x, I171x, I172x, I173x, I174x, I175x, I176x, I177x, I178x, I179x, I180x, I181x, I182x, I183x, I184x, I185x, I186x;
always@(posedge clk)
	begin
	I0x = 8'd61;
	I1x = 8'd60;
	I2x = 8'd41;
	I3x = 8'd19;
	I4x = 8'd4;
	I5x = 8'd0;
	I6x = 8'd3;
	I7x = 8'd6;
	I8x = 8'd6;
	I9x = 8'd6;
	I10x = 8'd6;
	I11x = 8'd6;
	I12x = 8'd7;
	I13x = 8'd7;
	I14x = 8'd7;
	I15x = 8'd8;
	I16x = 8'd8;
	I17x = 8'd8;
	I18x = 8'd8;
	I19x = 8'd8;
	I20x = 8'd9;
	I21x = 8'd10;
	I22x = 8'd10;
	I23x = 8'd11;
	I24x = 8'd11;
	I25x = 8'd12;
	I26x = 8'd13;
	I27x = 8'd14;
	I28x = 8'd15;
	I29x = 8'd17;
	I30x = 8'd18;
	I31x = 8'd20;
	I32x = 8'd21;
	I33x = 8'd22;
	I34x = 8'd23;
	I35x = 8'd23;
	I36x = 8'd23;
	I37x = 8'd22;
	I38x = 8'd21;
	I39x = 8'd19;
	I40x = 8'd16;
	I41x = 8'd14;
	I42x = 8'd12;
	I43x = 8'd11;
	I44x = 8'd9;
	I45x = 8'd9;
	I46x = 8'd8;
	I47x = 8'd7;
	I48x = 8'd7;
	I49x = 8'd7;
	I50x = 8'd7;
	I51x = 8'd7;
	I52x = 8'd7;
	I53x = 8'd7;
	I54x = 8'd7;
	I55x = 8'd7;
	I56x = 8'd7;
	I57x = 8'd7;
	I58x = 8'd7;
	I59x = 8'd7;
	I60x = 8'd7;
	I61x = 8'd7;
	I62x = 8'd7;
	I63x = 8'd7;
	I64x = 8'd7;
	I65x = 8'd7;
	I66x = 8'd7;
	I67x = 8'd7;
	I68x = 8'd7;
	I69x = 8'd7;
	I70x = 8'd7;
	I71x = 8'd6;
	I72x = 8'd7;
	I73x = 8'd6;
	I74x = 8'd6;
	I75x = 8'd6;
	I76x = 8'd6;
	I77x = 8'd6;
	I78x = 8'd6;
	I79x = 8'd6;
	I80x = 8'd6;
	I81x = 8'd6;
	I82x = 8'd6;
	I83x = 8'd6;
	I84x = 8'd6;
	I85x = 8'd6;
	I86x = 8'd6;
	I87x = 8'd6;
	I88x = 8'd6;
	I89x = 8'd6;
	I90x = 8'd6;
	I91x = 8'd6;
	I92x = 8'd6;
	I93x = 8'd6;
	I94x = 8'd6;
	I95x = 8'd6;
	I96x = 8'd6;
	I97x = 8'd6;
	I98x = 8'd6;
	I99x = 8'd6;
	I100x = 8'd6;
	I101x = 8'd6;
	I102x = 8'd6;
	I103x = 8'd6;
	I104x = 8'd6;
	I105x = 8'd6;
	I106x = 8'd7;
	I107x = 8'd8;
	I108x = 8'd10;
	I109x = 8'd11;
	I110x = 8'd12;
	I111x = 8'd14;
	I112x = 8'd15;
	I113x = 8'd14;
	I114x = 8'd14;
	I115x = 8'd12;
	I116x = 8'd11;
	I117x = 8'd10;
	I118x = 8'd7;
	I119x = 8'd6;
	I120x = 8'd5;
	I121x = 8'd5;
	I122x = 8'd5;
	I123x = 8'd5;
	I124x = 8'd5;
	I125x = 8'd3;
	I126x = 8'd5;
	I127x = 8'd17;
	I128x = 8'd46;
	I129x = 8'd64;
	I130x = 8'd58;
	I131x = 8'd31;
	I132x = 8'd14;
	I133x = 8'd2;
	I134x = 8'd3;
	I135x = 8'd7;
	I136x = 8'd8;
	I137x = 8'd7;
	I138x = 8'd8;
	I139x = 8'd8;
	I140x = 8'd8;
	I141x = 8'd8;
	I142x = 8'd9;
	I143x = 8'd9;
	I144x = 8'd9;
	I145x = 8'd10;
	I146x = 8'd10;
	I147x = 8'd10;
	I148x = 8'd11;
	I149x = 8'd11;
	I150x = 8'd12;
	I151x = 8'd12;
	I152x = 8'd13;
	I153x = 8'd14;
	I154x = 8'd0;
	I155x = 8'd0;
	I156x = 8'd0;
	I157x = 8'd0;
	I158x = 8'd0;
	I159x = 8'd0;
	I160x = 8'd0;
	I161x = 8'd0;
	I162x = 8'd0;
	I163x = 8'd0;
	I164x = 8'd0;
	I165x = 8'd0;
	I166x = 8'd0;
	I167x = 8'd0;
	I168x = 8'd0;
	I169x = 8'd0;
	I170x = 8'd0;
	I171x = 8'd0;
	I172x = 8'd0;
	I173x = 8'd0;
	I174x = 8'd0;
	I175x = 8'd0;
	I176x = 8'd0;
	I177x = 8'd0;
	I178x = 8'd0;
	I179x = 8'd0;
	I180x = 8'd0;
	I181x = 8'd0;
	I182x = 8'd0;
	I183x = 8'd0;
	I184x = 8'd0;
	I185x = 8'd0;
	I186x = 8'd0;
	end
endmodule
