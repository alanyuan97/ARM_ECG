module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = -6909;
	I1x = 1516;
	I2x = 3071;
	I3x = -3580;
	I4x = -2036;
	I5x = -1257;
	I6x = 3366;
	I7x = 6191;
	I8x = 3743;
	I9x = 8183;
	I10x = 2420;
	I11x = -3089;
	I12x = 6716;
	I13x = -6712;
	I14x = -6874;
	I15x = 1474;
	I16x = 775;
	I17x = 1943;
	I18x = 4393;
	I19x = -6397;
	I20x = -2688;
	I21x = 2177;
	I22x = 136;
	I23x = -5340;
	I24x = -4398;
	I25x = -6181;
	I26x = -4251;
	I27x = -6457;
	I28x = 2227;
	I29x = -6314;
	I30x = -6242;
	I31x = -2902;
	I32x = 4957;
	I33x = 6201;
	I34x = 4399;
	I35x = -6865;
	I36x = -4136;
	I37x = 7847;
	I38x = 8133;
	I39x = 1443;
	I40x = 445;
	I41x = -6253;
	I42x = -2923;
	I43x = -6443;
	I44x = 4800;
	I45x = 5899;
	I46x = -1408;
	I47x = -4729;
	I48x = 6354;
	I49x = -4920;
	I50x = -203;
	I51x = 1374;
	I52x = -7865;
	I53x = 7438;
	I54x = 2771;
	I55x = 6310;
	I56x = -1317;
	I57x = 3104;
	I58x = -7883;
	I59x = 3735;
	I60x = -6935;
	I61x = -7696;
	I62x = 7057;
	I63x = 4464;
	I64x = 5638;
	I65x = 140;
	I66x = 4922;
	I67x = 4175;
	I68x = 5289;
	I69x = -6139;
	I70x = -7586;
	I71x = -7095;
	I72x = -5087;
	I73x = 2207;
	I74x = -6804;
	I75x = 5247;
	I76x = -6177;
	I77x = 4007;
	I78x = -3262;
	I79x = -351;
	I80x = 7612;
	I81x = 7556;
	I82x = -4178;
	I83x = -7636;
	I84x = 2401;
	I85x = -2989;
	I86x = -1947;
	I87x = 8046;
	I88x = 2117;
	I89x = -5378;
	I90x = -1641;
	I91x = 6484;
	I92x = -5480;
	I93x = 4855;
	I94x = 3573;
	I95x = 4979;
	I96x = 4632;
	I97x = -4102;
	I98x = -4406;
	I99x = 6627;
	I100x = 5669;
	I101x = 6426;
	I102x = -7274;
	I103x = 4323;
	I104x = 794;
	I105x = -293;
	I106x = 7089;
	I107x = -545;
	I108x = 5129;
	I109x = -2786;
	I110x = -7083;
	I111x = 5636;
	I112x = -6678;
	I113x = -3787;
	I114x = 1717;
	I115x = -6942;
	I116x = 5394;
	I117x = 3961;
	I118x = 348;
	I119x = -5180;
	I120x = 1965;
	I121x = -562;
	I122x = -146;
	I123x = 928;
	I124x = -1606;
	I125x = 1837;
	I126x = 4900;
	I127x = -3166;
	I128x = 292;
	I129x = -7521;
	I130x = -3484;
	I131x = -1670;
	I132x = -4745;
	I133x = 5348;
	I134x = 4904;
	I135x = 6373;
	I136x = -3349;
	I137x = 7961;
	I138x = -1630;
	I139x = 7324;
	I140x = 443;
	I141x = -3624;
	I142x = 870;
	I143x = -4446;
	I144x = -7593;
	I145x = -8025;
	I146x = -1072;
	I147x = -383;
	I148x = -6006;
	I149x = -4282;
	I150x = 4800;
	I151x = 2562;
	I152x = -5491;
	I153x = -5455;
	I154x = 3830;
	I155x = 2183;
	I156x = 5978;
	I157x = 5332;
	I158x = 2709;
	I159x = -4412;
	I160x = 6482;
	I161x = 5316;
	I162x = -2799;
	I163x = 2925;
	I164x = -3878;
	I165x = 486;
	I166x = 2092;
	I167x = 5956;
	I168x = -3335;
	I169x = 2299;
	I170x = -7036;
	I171x = -5184;
	I172x = -7132;
	I173x = -5100;
	I174x = 8101;
	I175x = 2841;
	I176x = 2880;
	I177x = 1981;
	I178x = -7640;
	I179x = -5144;
	I180x = -1126;
	I181x = 5297;
	I182x = 1011;
	I183x = -1273;
	I184x = 3096;
	I185x = -3819;
	I186x = -5243;
	end
endmodule
[0.39406153 0.56610646 0.         0.         1.55277877] 

 [3228, 4637, 0, 0, 12720] 

 ['0000110010011100', '0001001000011101', '0000000000000000', '0000000000000000', '0011000110110000']
