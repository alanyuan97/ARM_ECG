module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 1004;
	I1x = 786;
	I2x = 394;
	I3x = 179;
	I4x = 0;
	I5x = 13;
	I6x = 74;
	I7x = 111;
	I8x = 118;
	I9x = 135;
	I10x = 142;
	I11x = 146;
	I12x = 154;
	I13x = 154;
	I14x = 149;
	I15x = 161;
	I16x = 167;
	I17x = 176;
	I18x = 181;
	I19x = 189;
	I20x = 195;
	I21x = 206;
	I22x = 219;
	I23x = 227;
	I24x = 256;
	I25x = 280;
	I26x = 303;
	I27x = 324;
	I28x = 359;
	I29x = 366;
	I30x = 390;
	I31x = 411;
	I32x = 427;
	I33x = 428;
	I34x = 417;
	I35x = 413;
	I36x = 382;
	I37x = 347;
	I38x = 309;
	I39x = 275;
	I40x = 243;
	I41x = 235;
	I42x = 215;
	I43x = 198;
	I44x = 198;
	I45x = 188;
	I46x = 181;
	I47x = 176;
	I48x = 179;
	I49x = 176;
	I50x = 177;
	I51x = 177;
	I52x = 192;
	I53x = 198;
	I54x = 188;
	I55x = 187;
	I56x = 182;
	I57x = 188;
	I58x = 195;
	I59x = 194;
	I60x = 190;
	I61x = 181;
	I62x = 186;
	I63x = 175;
	I64x = 185;
	I65x = 188;
	I66x = 181;
	I67x = 173;
	I68x = 181;
	I69x = 190;
	I70x = 185;
	I71x = 185;
	I72x = 189;
	I73x = 190;
	I74x = 196;
	I75x = 192;
	I76x = 192;
	I77x = 196;
	I78x = 191;
	I79x = 192;
	I80x = 184;
	I81x = 201;
	I82x = 215;
	I83x = 232;
	I84x = 253;
	I85x = 284;
	I86x = 305;
	I87x = 328;
	I88x = 321;
	I89x = 321;
	I90x = 277;
	I91x = 263;
	I92x = 242;
	I93x = 196;
	I94x = 163;
	I95x = 158;
	I96x = 161;
	I97x = 154;
	I98x = 162;
	I99x = 154;
	I100x = 148;
	I101x = 118;
	I102x = 163;
	I103x = 424;
	I104x = 867;
	I105x = 1024;
	I106x = 785;
	I107x = 419;
	I108x = 222;
	I109x = 42;
	I110x = 54;
	I111x = 120;
	I112x = 155;
	I113x = 160;
	I114x = 163;
	I115x = 166;
	I116x = 176;
	I117x = 178;
	I118x = 184;
	I119x = 185;
	I120x = 182;
	I121x = 179;
	I122x = 195;
	I123x = 195;
	I124x = 208;
	I125x = 208;
	I126x = 220;
	I127x = 236;
	I128x = 244;
	I129x = 257;
	I130x = 272;
	I131x = 296;
	I132x = 318;
	I133x = 338;
	I134x = 368;
	I135x = 385;
	I136x = 399;
	I137x = 409;
	I138x = 414;
	I139x = 416;
	I140x = 401;
	I141x = 378;
	I142x = 348;
	I143x = 318;
	I144x = 0;
	I145x = 0;
	I146x = 0;
	I147x = 0;
	I148x = 0;
	I149x = 0;
	I150x = 0;
	I151x = 0;
	I152x = 0;
	I153x = 0;
	I154x = 0;
	I155x = 0;
	I156x = 0;
	I157x = 0;
	I158x = 0;
	I159x = 0;
	I160x = 0;
	I161x = 0;
	I162x = 0;
	I163x = 0;
	I164x = 0;
	I165x = 0;
	I166x = 0;
	I167x = 0;
	I168x = 0;
	I169x = 0;
	I170x = 0;
	I171x = 0;
	I172x = 0;
	I173x = 0;
	I174x = 0;
	I175x = 0;
	I176x = 0;
	I177x = 0;
	I178x = 0;
	I179x = 0;
	I180x = 0;
	I181x = 0;
	I182x = 0;
	I183x = 0;
	I184x = 0;
	I185x = 0;
	I186x = 0;
	end
endmodule
