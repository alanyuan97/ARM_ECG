module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x);
	input EN;
	output reg [23:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x;
	always@(negedge EN)
		begin
			   I0x <= 22;      //expecting 1
				I1x <= 8;
				I2x <= -1;
				I3x <= 6;
				I4x <= 3;
				I5x <= 6;
				I6x <= 4;
				I7x <= 6;
				I8x <= 5;
				I9x <= 7;
				I10x <= 6;
				I11x <= 8;
				I12x <= 9;
				I13x <= 13;
				I14x <= 14;
				I15x <= 16;
				I16x <= 12;
				I17x <= 9;
				I18x <= 5;
				I19x <= 4;
				I20x <= 3;
				I21x <= 3;
				I22x <= 3;
				I23x <= 4;
				I24x <= 3;
				I25x <= 4;
				I26x <= 3;
				I27x <= 4;
				I28x <= 3;
				I29x <= 3;
				I30x <= 2;
				I31x <= 3;
				I32x <= 2;
				I33x <= 2;
				I34x <= 2;
				I35x <= 3;
				I36x <= 2;
				I37x <= 3;
				I38x <= 2;
				I39x <= 3;
				I40x <= 2;
				I41x <= 3;
				I42x <= 4;
				I43x <= 6;
				I44x <= 5;
				I45x <= 4;
				I46x <= 2;
				I47x <= 3;
				I48x <= 2;
				I49x <= 3;
				I50x <= 1;
				I51x <= 27;
				I52x <= 6;
				I53x <= 0;
				I54x <= 6;
				I55x <= 4;
				I56x <= 5;
				I57x <= 5;
				I58x <= 6;
				I59x <= 6;
				I60x <= 7;
				I61x <= 2;
				I62x <= 0;
				I63x <= 0;
				I64x <= 0;
				I65x <= 0;
				I66x <= 0;
				I67x <= 0;
				I68x <= 0;
				I69x <= 0;
				I70x <= 0;
				I71x <= 0;
				I72x <= -1;
				I73x <= 1;
				I74x <= -2;
	end
endmodule
