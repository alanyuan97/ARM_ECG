module node_1_3(clk,reset,N3x,A0x,A1x,A2x,A3x,A4x,A5x,A6x,A7x,A8x,A9x,A10x,A11x,A12x,A13x,A14x,A15x,A16x,A17x,A18x,A19x,A20x,A21x,A22x,A23x,A24x,A25x,A26x,A27x,A28x,A29x,A30x,A31x,A32x,A33x,A34x,A35x,A36x,A37x,A38x,A39x,A40x,A41x,A42x,A43x,A44x,A45x,A46x,A47x,A48x,A49x,A50x,A51x,A52x,A53x,A54x,A55x,A56x,A57x,A58x,A59x,A60x,A61x,A62x,A63x,A64x,A65x,A66x,A67x,A68x,A69x,A70x,A71x,A72x,A73x,A74x,A75x,A76x,A77x,A78x,A79x,A80x,A81x,A82x,A83x,A84x,A85x,A86x,A87x,A88x,A89x,A90x,A91x,A92x,A93x,A94x,A95x,A96x,A97x,A98x,A99x,A100x,A101x,A102x,A103x,A104x,A105x,A106x,A107x,A108x,A109x,A110x,A111x,A112x,A113x,A114x,A115x,A116x,A117x,A118x,A119x,A120x,A121x,A122x,A123x,A124x,A125x,A126x,A127x,A128x,A129x,A130x,A131x,A132x,A133x,A134x,A135x,A136x,A137x,A138x,A139x,A140x,A141x,A142x,A143x,A144x,A145x,A146x,A147x,A148x,A149x,A150x,A151x,A152x,A153x,A154x,A155x,A156x,A157x,A158x,A159x,A160x,A161x,A162x,A163x,A164x,A165x,A166x,A167x,A168x,A169x,A170x,A171x,A172x,A173x,A174x,A175x,A176x,A177x,A178x,A179x,A180x,A181x,A182x,A183x,A184x,A185x,A186x);
	input clk;
	input reset;
	input [7:0] A0x, A1x, A2x, A3x, A4x, A5x, A6x, A7x, A8x, A9x, A10x, A11x, A12x, A13x, A14x, A15x, A16x, A17x, A18x, A19x, A20x, A21x, A22x, A23x, A24x, A25x, A26x, A27x, A28x, A29x, A30x, A31x, A32x, A33x, A34x, A35x, A36x, A37x, A38x, A39x, A40x, A41x, A42x, A43x, A44x, A45x, A46x, A47x, A48x, A49x, A50x, A51x, A52x, A53x, A54x, A55x, A56x, A57x, A58x, A59x, A60x, A61x, A62x, A63x, A64x, A65x, A66x, A67x, A68x, A69x, A70x, A71x, A72x, A73x, A74x, A75x, A76x, A77x, A78x, A79x, A80x, A81x, A82x, A83x, A84x, A85x, A86x, A87x, A88x, A89x, A90x, A91x, A92x, A93x, A94x, A95x, A96x, A97x, A98x, A99x, A100x, A101x, A102x, A103x, A104x, A105x, A106x, A107x, A108x, A109x, A110x, A111x, A112x, A113x, A114x, A115x, A116x, A117x, A118x, A119x, A120x, A121x, A122x, A123x, A124x, A125x, A126x, A127x, A128x, A129x, A130x, A131x, A132x, A133x, A134x, A135x, A136x, A137x, A138x, A139x, A140x, A141x, A142x, A143x, A144x, A145x, A146x, A147x, A148x, A149x, A150x, A151x, A152x, A153x, A154x, A155x, A156x, A157x, A158x, A159x, A160x, A161x, A162x, A163x, A164x, A165x, A166x, A167x, A168x, A169x, A170x, A171x, A172x, A173x, A174x, A175x, A176x, A177x, A178x, A179x, A180x, A181x, A182x, A183x, A184x, A185x, A186x;
	reg [7:0] A0x_c, A1x_c, A2x_c, A3x_c, A4x_c, A5x_c, A6x_c, A7x_c, A8x_c, A9x_c, A10x_c, A11x_c, A12x_c, A13x_c, A14x_c, A15x_c, A16x_c, A17x_c, A18x_c, A19x_c, A20x_c, A21x_c, A22x_c, A23x_c, A24x_c, A25x_c, A26x_c, A27x_c, A28x_c, A29x_c, A30x_c, A31x_c, A32x_c, A33x_c, A34x_c, A35x_c, A36x_c, A37x_c, A38x_c, A39x_c, A40x_c, A41x_c, A42x_c, A43x_c, A44x_c, A45x_c, A46x_c, A47x_c, A48x_c, A49x_c, A50x_c, A51x_c, A52x_c, A53x_c, A54x_c, A55x_c, A56x_c, A57x_c, A58x_c, A59x_c, A60x_c, A61x_c, A62x_c, A63x_c, A64x_c, A65x_c, A66x_c, A67x_c, A68x_c, A69x_c, A70x_c, A71x_c, A72x_c, A73x_c, A74x_c, A75x_c, A76x_c, A77x_c, A78x_c, A79x_c, A80x_c, A81x_c, A82x_c, A83x_c, A84x_c, A85x_c, A86x_c, A87x_c, A88x_c, A89x_c, A90x_c, A91x_c, A92x_c, A93x_c, A94x_c, A95x_c, A96x_c, A97x_c, A98x_c, A99x_c, A100x_c, A101x_c, A102x_c, A103x_c, A104x_c, A105x_c, A106x_c, A107x_c, A108x_c, A109x_c, A110x_c, A111x_c, A112x_c, A113x_c, A114x_c, A115x_c, A116x_c, A117x_c, A118x_c, A119x_c, A120x_c, A121x_c, A122x_c, A123x_c, A124x_c, A125x_c, A126x_c, A127x_c, A128x_c, A129x_c, A130x_c, A131x_c, A132x_c, A133x_c, A134x_c, A135x_c, A136x_c, A137x_c, A138x_c, A139x_c, A140x_c, A141x_c, A142x_c, A143x_c, A144x_c, A145x_c, A146x_c, A147x_c, A148x_c, A149x_c, A150x_c, A151x_c, A152x_c, A153x_c, A154x_c, A155x_c, A156x_c, A157x_c, A158x_c, A159x_c, A160x_c, A161x_c, A162x_c, A163x_c, A164x_c, A165x_c, A166x_c, A167x_c, A168x_c, A169x_c, A170x_c, A171x_c, A172x_c, A173x_c, A174x_c, A175x_c, A176x_c, A177x_c, A178x_c, A179x_c, A180x_c, A181x_c, A182x_c, A183x_c, A184x_c, A185x_c, A186x_c;
	wire [15:0] sum0x, sum1x, sum2x, sum3x, sum4x, sum5x, sum6x, sum7x, sum8x, sum9x, sum10x, sum11x, sum12x, sum13x, sum14x, sum15x, sum16x, sum17x, sum18x, sum19x, sum20x, sum21x, sum22x, sum23x, sum24x, sum25x, sum26x, sum27x, sum28x, sum29x, sum30x, sum31x, sum32x, sum33x, sum34x, sum35x, sum36x, sum37x, sum38x, sum39x, sum40x, sum41x, sum42x, sum43x, sum44x, sum45x, sum46x, sum47x, sum48x, sum49x, sum50x, sum51x, sum52x, sum53x, sum54x, sum55x, sum56x, sum57x, sum58x, sum59x, sum60x, sum61x, sum62x, sum63x, sum64x, sum65x, sum66x, sum67x, sum68x, sum69x, sum70x, sum71x, sum72x, sum73x, sum74x, sum75x, sum76x, sum77x, sum78x, sum79x, sum80x, sum81x, sum82x, sum83x, sum84x, sum85x, sum86x, sum87x, sum88x, sum89x, sum90x, sum91x, sum92x, sum93x, sum94x, sum95x, sum96x, sum97x, sum98x, sum99x, sum100x, sum101x, sum102x, sum103x, sum104x, sum105x, sum106x, sum107x, sum108x, sum109x, sum110x, sum111x, sum112x, sum113x, sum114x, sum115x, sum116x, sum117x, sum118x, sum119x, sum120x, sum121x, sum122x, sum123x, sum124x, sum125x, sum126x, sum127x, sum128x, sum129x, sum130x, sum131x, sum132x, sum133x, sum134x, sum135x, sum136x, sum137x, sum138x, sum139x, sum140x, sum141x, sum142x, sum143x, sum144x, sum145x, sum146x, sum147x, sum148x, sum149x, sum150x, sum151x, sum152x, sum153x, sum154x, sum155x, sum156x, sum157x, sum158x, sum159x, sum160x, sum161x, sum162x, sum163x, sum164x, sum165x, sum166x, sum167x, sum168x, sum169x, sum170x, sum171x, sum172x, sum173x, sum174x, sum175x, sum176x, sum177x, sum178x, sum179x, sum180x, sum181x, sum182x, sum183x, sum184x, sum185x, sum186x;
	output reg [7:0] N3x;
	reg [22:0] sumout;

	parameter [7:0] W0x=-8'd11;
	parameter [7:0] W1x=-8'd31;
	parameter [7:0] W2x=8'd19;
	parameter [7:0] W3x=8'd25;
	parameter [7:0] W4x=8'd27;
	parameter [7:0] W5x=8'd18;
	parameter [7:0] W6x=-8'd1;
	parameter [7:0] W7x=-8'd16;
	parameter [7:0] W8x=8'd2;
	parameter [7:0] W9x=-8'd11;
	parameter [7:0] W10x=-8'd14;
	parameter [7:0] W11x=-8'd13;
	parameter [7:0] W12x=-8'd13;
	parameter [7:0] W13x=-8'd9;
	parameter [7:0] W14x=-8'd7;
	parameter [7:0] W15x=-8'd2;
	parameter [7:0] W16x=8'd3;
	parameter [7:0] W17x=-8'd10;
	parameter [7:0] W18x=-8'd5;
	parameter [7:0] W19x=8'd0;
	parameter [7:0] W20x=8'd9;
	parameter [7:0] W21x=8'd5;
	parameter [7:0] W22x=8'd12;
	parameter [7:0] W23x=-8'd5;
	parameter [7:0] W24x=-8'd5;
	parameter [7:0] W25x=8'd10;
	parameter [7:0] W26x=8'd9;
	parameter [7:0] W27x=8'd7;
	parameter [7:0] W28x=8'd12;
	parameter [7:0] W29x=8'd11;
	parameter [7:0] W30x=8'd10;
	parameter [7:0] W31x=8'd12;
	parameter [7:0] W32x=8'd2;
	parameter [7:0] W33x=8'd10;
	parameter [7:0] W34x=8'd14;
	parameter [7:0] W35x=8'd24;
	parameter [7:0] W36x=8'd17;
	parameter [7:0] W37x=8'd12;
	parameter [7:0] W38x=8'd7;
	parameter [7:0] W39x=8'd8;
	parameter [7:0] W40x=8'd13;
	parameter [7:0] W41x=8'd2;
	parameter [7:0] W42x=8'd9;
	parameter [7:0] W43x=-8'd6;
	parameter [7:0] W44x=8'd12;
	parameter [7:0] W45x=8'd10;
	parameter [7:0] W46x=8'd8;
	parameter [7:0] W47x=8'd11;
	parameter [7:0] W48x=8'd12;
	parameter [7:0] W49x=8'd4;
	parameter [7:0] W50x=8'd9;
	parameter [7:0] W51x=8'd10;
	parameter [7:0] W52x=8'd7;
	parameter [7:0] W53x=8'd11;
	parameter [7:0] W54x=-8'd6;
	parameter [7:0] W55x=-8'd11;
	parameter [7:0] W56x=8'd1;
	parameter [7:0] W57x=-8'd6;
	parameter [7:0] W58x=-8'd6;
	parameter [7:0] W59x=-8'd4;
	parameter [7:0] W60x=-8'd11;
	parameter [7:0] W61x=-8'd5;
	parameter [7:0] W62x=-8'd5;
	parameter [7:0] W63x=-8'd9;
	parameter [7:0] W64x=-8'd9;
	parameter [7:0] W65x=-8'd1;
	parameter [7:0] W66x=-8'd7;
	parameter [7:0] W67x=8'd7;
	parameter [7:0] W68x=8'd3;
	parameter [7:0] W69x=8'd6;
	parameter [7:0] W70x=8'd9;
	parameter [7:0] W71x=8'd13;
	parameter [7:0] W72x=-8'd4;
	parameter [7:0] W73x=-8'd2;
	parameter [7:0] W74x=8'd6;
	parameter [7:0] W75x=8'd1;
	parameter [7:0] W76x=-8'd1;
	parameter [7:0] W77x=8'd6;
	parameter [7:0] W78x=8'd6;
	parameter [7:0] W79x=8'd2;
	parameter [7:0] W80x=8'd7;
	parameter [7:0] W81x=8'd2;
	parameter [7:0] W82x=8'd7;
	parameter [7:0] W83x=8'd2;
	parameter [7:0] W84x=8'd10;
	parameter [7:0] W85x=-8'd2;
	parameter [7:0] W86x=-8'd18;
	parameter [7:0] W87x=-8'd5;
	parameter [7:0] W88x=8'd0;
	parameter [7:0] W89x=-8'd9;
	parameter [7:0] W90x=8'd2;
	parameter [7:0] W91x=-8'd4;
	parameter [7:0] W92x=8'd0;
	parameter [7:0] W93x=8'd0;
	parameter [7:0] W94x=8'd7;
	parameter [7:0] W95x=8'd0;
	parameter [7:0] W96x=-8'd1;
	parameter [7:0] W97x=8'd9;
	parameter [7:0] W98x=8'd4;
	parameter [7:0] W99x=8'd2;
	parameter [7:0] W100x=8'd3;
	parameter [7:0] W101x=8'd3;
	parameter [7:0] W102x=8'd8;
	parameter [7:0] W103x=8'd3;
	parameter [7:0] W104x=8'd12;
	parameter [7:0] W105x=8'd0;
	parameter [7:0] W106x=8'd18;
	parameter [7:0] W107x=8'd2;
	parameter [7:0] W108x=-8'd6;
	parameter [7:0] W109x=8'd8;
	parameter [7:0] W110x=-8'd2;
	parameter [7:0] W111x=-8'd5;
	parameter [7:0] W112x=-8'd4;
	parameter [7:0] W113x=-8'd5;
	parameter [7:0] W114x=-8'd17;
	parameter [7:0] W115x=-8'd7;
	parameter [7:0] W116x=-8'd5;
	parameter [7:0] W117x=-8'd3;
	parameter [7:0] W118x=8'd0;
	parameter [7:0] W119x=8'd3;
	parameter [7:0] W120x=8'd6;
	parameter [7:0] W121x=-8'd4;
	parameter [7:0] W122x=8'd8;
	parameter [7:0] W123x=8'd5;
	parameter [7:0] W124x=-8'd9;
	parameter [7:0] W125x=8'd9;
	parameter [7:0] W126x=-8'd5;
	parameter [7:0] W127x=8'd6;
	parameter [7:0] W128x=-8'd1;
	parameter [7:0] W129x=8'd0;
	parameter [7:0] W130x=8'd7;
	parameter [7:0] W131x=-8'd6;
	parameter [7:0] W132x=-8'd4;
	parameter [7:0] W133x=8'd3;
	parameter [7:0] W134x=8'd7;
	parameter [7:0] W135x=-8'd9;
	parameter [7:0] W136x=8'd6;
	parameter [7:0] W137x=-8'd2;
	parameter [7:0] W138x=8'd12;
	parameter [7:0] W139x=-8'd4;
	parameter [7:0] W140x=-8'd3;
	parameter [7:0] W141x=-8'd5;
	parameter [7:0] W142x=8'd11;
	parameter [7:0] W143x=-8'd6;
	parameter [7:0] W144x=8'd11;
	parameter [7:0] W145x=-8'd2;
	parameter [7:0] W146x=8'd8;
	parameter [7:0] W147x=8'd8;
	parameter [7:0] W148x=8'd20;
	parameter [7:0] W149x=8'd5;
	parameter [7:0] W150x=-8'd20;
	parameter [7:0] W151x=8'd3;
	parameter [7:0] W152x=-8'd7;
	parameter [7:0] W153x=-8'd15;
	parameter [7:0] W154x=-8'd5;
	parameter [7:0] W155x=-8'd16;
	parameter [7:0] W156x=8'd7;
	parameter [7:0] W157x=-8'd31;
	parameter [7:0] W158x=-8'd31;
	parameter [7:0] W159x=-8'd20;
	parameter [7:0] W160x=-8'd6;
	parameter [7:0] W161x=-8'd7;
	parameter [7:0] W162x=-8'd8;
	parameter [7:0] W163x=-8'd24;
	parameter [7:0] W164x=-8'd10;
	parameter [7:0] W165x=-8'd6;
	parameter [7:0] W166x=-8'd4;
	parameter [7:0] W167x=8'd7;
	parameter [7:0] W168x=8'd0;
	parameter [7:0] W169x=8'd7;
	parameter [7:0] W170x=-8'd13;
	parameter [7:0] W171x=8'd3;
	parameter [7:0] W172x=8'd14;
	parameter [7:0] W173x=8'd9;
	parameter [7:0] W174x=8'd2;
	parameter [7:0] W175x=-8'd8;
	parameter [7:0] W176x=-8'd12;
	parameter [7:0] W177x=-8'd29;
	parameter [7:0] W178x=-8'd25;
	parameter [7:0] W179x=-8'd11;
	parameter [7:0] W180x=-8'd24;
	parameter [7:0] W181x=-8'd9;
	parameter [7:0] W182x=-8'd18;
	parameter [7:0] W183x=-8'd18;
	parameter [7:0] W184x=-8'd14;
	parameter [7:0] W185x=-8'd15;
	parameter [7:0] W186x=-8'd11;
	parameter [15:0] B0x=-16'd1024;


	assign sum0x = {A0x_c[7],A0x_c[7],A0x_c[7],A0x_c[7],A0x_c[7],A0x_c[7],A0x_c[7],A0x_c[7],A0x_c}*{W0x[7],W0x[7],W0x[7],W0x[7],W0x[7],W0x[7],W0x[7],W0x[7],W0x};
	assign sum1x = {A1x_c[7],A1x_c[7],A1x_c[7],A1x_c[7],A1x_c[7],A1x_c[7],A1x_c[7],A1x_c[7],A1x_c}*{W1x[7],W1x[7],W1x[7],W1x[7],W1x[7],W1x[7],W1x[7],W1x[7],W1x};
	assign sum2x = {A2x_c[7],A2x_c[7],A2x_c[7],A2x_c[7],A2x_c[7],A2x_c[7],A2x_c[7],A2x_c[7],A2x_c}*{W2x[7],W2x[7],W2x[7],W2x[7],W2x[7],W2x[7],W2x[7],W2x[7],W2x};
	assign sum3x = {A3x_c[7],A3x_c[7],A3x_c[7],A3x_c[7],A3x_c[7],A3x_c[7],A3x_c[7],A3x_c[7],A3x_c}*{W3x[7],W3x[7],W3x[7],W3x[7],W3x[7],W3x[7],W3x[7],W3x[7],W3x};
	assign sum4x = {A4x_c[7],A4x_c[7],A4x_c[7],A4x_c[7],A4x_c[7],A4x_c[7],A4x_c[7],A4x_c[7],A4x_c}*{W4x[7],W4x[7],W4x[7],W4x[7],W4x[7],W4x[7],W4x[7],W4x[7],W4x};
	assign sum5x = {A5x_c[7],A5x_c[7],A5x_c[7],A5x_c[7],A5x_c[7],A5x_c[7],A5x_c[7],A5x_c[7],A5x_c}*{W5x[7],W5x[7],W5x[7],W5x[7],W5x[7],W5x[7],W5x[7],W5x[7],W5x};
	assign sum6x = {A6x_c[7],A6x_c[7],A6x_c[7],A6x_c[7],A6x_c[7],A6x_c[7],A6x_c[7],A6x_c[7],A6x_c}*{W6x[7],W6x[7],W6x[7],W6x[7],W6x[7],W6x[7],W6x[7],W6x[7],W6x};
	assign sum7x = {A7x_c[7],A7x_c[7],A7x_c[7],A7x_c[7],A7x_c[7],A7x_c[7],A7x_c[7],A7x_c[7],A7x_c}*{W7x[7],W7x[7],W7x[7],W7x[7],W7x[7],W7x[7],W7x[7],W7x[7],W7x};
	assign sum8x = {A8x_c[7],A8x_c[7],A8x_c[7],A8x_c[7],A8x_c[7],A8x_c[7],A8x_c[7],A8x_c[7],A8x_c}*{W8x[7],W8x[7],W8x[7],W8x[7],W8x[7],W8x[7],W8x[7],W8x[7],W8x};
	assign sum9x = {A9x_c[7],A9x_c[7],A9x_c[7],A9x_c[7],A9x_c[7],A9x_c[7],A9x_c[7],A9x_c[7],A9x_c}*{W9x[7],W9x[7],W9x[7],W9x[7],W9x[7],W9x[7],W9x[7],W9x[7],W9x};
	assign sum10x = {A10x_c[7],A10x_c[7],A10x_c[7],A10x_c[7],A10x_c[7],A10x_c[7],A10x_c[7],A10x_c[7],A10x_c}*{W10x[7],W10x[7],W10x[7],W10x[7],W10x[7],W10x[7],W10x[7],W10x[7],W10x};
	assign sum11x = {A11x_c[7],A11x_c[7],A11x_c[7],A11x_c[7],A11x_c[7],A11x_c[7],A11x_c[7],A11x_c[7],A11x_c}*{W11x[7],W11x[7],W11x[7],W11x[7],W11x[7],W11x[7],W11x[7],W11x[7],W11x};
	assign sum12x = {A12x_c[7],A12x_c[7],A12x_c[7],A12x_c[7],A12x_c[7],A12x_c[7],A12x_c[7],A12x_c[7],A12x_c}*{W12x[7],W12x[7],W12x[7],W12x[7],W12x[7],W12x[7],W12x[7],W12x[7],W12x};
	assign sum13x = {A13x_c[7],A13x_c[7],A13x_c[7],A13x_c[7],A13x_c[7],A13x_c[7],A13x_c[7],A13x_c[7],A13x_c}*{W13x[7],W13x[7],W13x[7],W13x[7],W13x[7],W13x[7],W13x[7],W13x[7],W13x};
	assign sum14x = {A14x_c[7],A14x_c[7],A14x_c[7],A14x_c[7],A14x_c[7],A14x_c[7],A14x_c[7],A14x_c[7],A14x_c}*{W14x[7],W14x[7],W14x[7],W14x[7],W14x[7],W14x[7],W14x[7],W14x[7],W14x};
	assign sum15x = {A15x_c[7],A15x_c[7],A15x_c[7],A15x_c[7],A15x_c[7],A15x_c[7],A15x_c[7],A15x_c[7],A15x_c}*{W15x[7],W15x[7],W15x[7],W15x[7],W15x[7],W15x[7],W15x[7],W15x[7],W15x};
	assign sum16x = {A16x_c[7],A16x_c[7],A16x_c[7],A16x_c[7],A16x_c[7],A16x_c[7],A16x_c[7],A16x_c[7],A16x_c}*{W16x[7],W16x[7],W16x[7],W16x[7],W16x[7],W16x[7],W16x[7],W16x[7],W16x};
	assign sum17x = {A17x_c[7],A17x_c[7],A17x_c[7],A17x_c[7],A17x_c[7],A17x_c[7],A17x_c[7],A17x_c[7],A17x_c}*{W17x[7],W17x[7],W17x[7],W17x[7],W17x[7],W17x[7],W17x[7],W17x[7],W17x};
	assign sum18x = {A18x_c[7],A18x_c[7],A18x_c[7],A18x_c[7],A18x_c[7],A18x_c[7],A18x_c[7],A18x_c[7],A18x_c}*{W18x[7],W18x[7],W18x[7],W18x[7],W18x[7],W18x[7],W18x[7],W18x[7],W18x};
	assign sum19x = {A19x_c[7],A19x_c[7],A19x_c[7],A19x_c[7],A19x_c[7],A19x_c[7],A19x_c[7],A19x_c[7],A19x_c}*{W19x[7],W19x[7],W19x[7],W19x[7],W19x[7],W19x[7],W19x[7],W19x[7],W19x};
	assign sum20x = {A20x_c[7],A20x_c[7],A20x_c[7],A20x_c[7],A20x_c[7],A20x_c[7],A20x_c[7],A20x_c[7],A20x_c}*{W20x[7],W20x[7],W20x[7],W20x[7],W20x[7],W20x[7],W20x[7],W20x[7],W20x};
	assign sum21x = {A21x_c[7],A21x_c[7],A21x_c[7],A21x_c[7],A21x_c[7],A21x_c[7],A21x_c[7],A21x_c[7],A21x_c}*{W21x[7],W21x[7],W21x[7],W21x[7],W21x[7],W21x[7],W21x[7],W21x[7],W21x};
	assign sum22x = {A22x_c[7],A22x_c[7],A22x_c[7],A22x_c[7],A22x_c[7],A22x_c[7],A22x_c[7],A22x_c[7],A22x_c}*{W22x[7],W22x[7],W22x[7],W22x[7],W22x[7],W22x[7],W22x[7],W22x[7],W22x};
	assign sum23x = {A23x_c[7],A23x_c[7],A23x_c[7],A23x_c[7],A23x_c[7],A23x_c[7],A23x_c[7],A23x_c[7],A23x_c}*{W23x[7],W23x[7],W23x[7],W23x[7],W23x[7],W23x[7],W23x[7],W23x[7],W23x};
	assign sum24x = {A24x_c[7],A24x_c[7],A24x_c[7],A24x_c[7],A24x_c[7],A24x_c[7],A24x_c[7],A24x_c[7],A24x_c}*{W24x[7],W24x[7],W24x[7],W24x[7],W24x[7],W24x[7],W24x[7],W24x[7],W24x};
	assign sum25x = {A25x_c[7],A25x_c[7],A25x_c[7],A25x_c[7],A25x_c[7],A25x_c[7],A25x_c[7],A25x_c[7],A25x_c}*{W25x[7],W25x[7],W25x[7],W25x[7],W25x[7],W25x[7],W25x[7],W25x[7],W25x};
	assign sum26x = {A26x_c[7],A26x_c[7],A26x_c[7],A26x_c[7],A26x_c[7],A26x_c[7],A26x_c[7],A26x_c[7],A26x_c}*{W26x[7],W26x[7],W26x[7],W26x[7],W26x[7],W26x[7],W26x[7],W26x[7],W26x};
	assign sum27x = {A27x_c[7],A27x_c[7],A27x_c[7],A27x_c[7],A27x_c[7],A27x_c[7],A27x_c[7],A27x_c[7],A27x_c}*{W27x[7],W27x[7],W27x[7],W27x[7],W27x[7],W27x[7],W27x[7],W27x[7],W27x};
	assign sum28x = {A28x_c[7],A28x_c[7],A28x_c[7],A28x_c[7],A28x_c[7],A28x_c[7],A28x_c[7],A28x_c[7],A28x_c}*{W28x[7],W28x[7],W28x[7],W28x[7],W28x[7],W28x[7],W28x[7],W28x[7],W28x};
	assign sum29x = {A29x_c[7],A29x_c[7],A29x_c[7],A29x_c[7],A29x_c[7],A29x_c[7],A29x_c[7],A29x_c[7],A29x_c}*{W29x[7],W29x[7],W29x[7],W29x[7],W29x[7],W29x[7],W29x[7],W29x[7],W29x};
	assign sum30x = {A30x_c[7],A30x_c[7],A30x_c[7],A30x_c[7],A30x_c[7],A30x_c[7],A30x_c[7],A30x_c[7],A30x_c}*{W30x[7],W30x[7],W30x[7],W30x[7],W30x[7],W30x[7],W30x[7],W30x[7],W30x};
	assign sum31x = {A31x_c[7],A31x_c[7],A31x_c[7],A31x_c[7],A31x_c[7],A31x_c[7],A31x_c[7],A31x_c[7],A31x_c}*{W31x[7],W31x[7],W31x[7],W31x[7],W31x[7],W31x[7],W31x[7],W31x[7],W31x};
	assign sum32x = {A32x_c[7],A32x_c[7],A32x_c[7],A32x_c[7],A32x_c[7],A32x_c[7],A32x_c[7],A32x_c[7],A32x_c}*{W32x[7],W32x[7],W32x[7],W32x[7],W32x[7],W32x[7],W32x[7],W32x[7],W32x};
	assign sum33x = {A33x_c[7],A33x_c[7],A33x_c[7],A33x_c[7],A33x_c[7],A33x_c[7],A33x_c[7],A33x_c[7],A33x_c}*{W33x[7],W33x[7],W33x[7],W33x[7],W33x[7],W33x[7],W33x[7],W33x[7],W33x};
	assign sum34x = {A34x_c[7],A34x_c[7],A34x_c[7],A34x_c[7],A34x_c[7],A34x_c[7],A34x_c[7],A34x_c[7],A34x_c}*{W34x[7],W34x[7],W34x[7],W34x[7],W34x[7],W34x[7],W34x[7],W34x[7],W34x};
	assign sum35x = {A35x_c[7],A35x_c[7],A35x_c[7],A35x_c[7],A35x_c[7],A35x_c[7],A35x_c[7],A35x_c[7],A35x_c}*{W35x[7],W35x[7],W35x[7],W35x[7],W35x[7],W35x[7],W35x[7],W35x[7],W35x};
	assign sum36x = {A36x_c[7],A36x_c[7],A36x_c[7],A36x_c[7],A36x_c[7],A36x_c[7],A36x_c[7],A36x_c[7],A36x_c}*{W36x[7],W36x[7],W36x[7],W36x[7],W36x[7],W36x[7],W36x[7],W36x[7],W36x};
	assign sum37x = {A37x_c[7],A37x_c[7],A37x_c[7],A37x_c[7],A37x_c[7],A37x_c[7],A37x_c[7],A37x_c[7],A37x_c}*{W37x[7],W37x[7],W37x[7],W37x[7],W37x[7],W37x[7],W37x[7],W37x[7],W37x};
	assign sum38x = {A38x_c[7],A38x_c[7],A38x_c[7],A38x_c[7],A38x_c[7],A38x_c[7],A38x_c[7],A38x_c[7],A38x_c}*{W38x[7],W38x[7],W38x[7],W38x[7],W38x[7],W38x[7],W38x[7],W38x[7],W38x};
	assign sum39x = {A39x_c[7],A39x_c[7],A39x_c[7],A39x_c[7],A39x_c[7],A39x_c[7],A39x_c[7],A39x_c[7],A39x_c}*{W39x[7],W39x[7],W39x[7],W39x[7],W39x[7],W39x[7],W39x[7],W39x[7],W39x};
	assign sum40x = {A40x_c[7],A40x_c[7],A40x_c[7],A40x_c[7],A40x_c[7],A40x_c[7],A40x_c[7],A40x_c[7],A40x_c}*{W40x[7],W40x[7],W40x[7],W40x[7],W40x[7],W40x[7],W40x[7],W40x[7],W40x};
	assign sum41x = {A41x_c[7],A41x_c[7],A41x_c[7],A41x_c[7],A41x_c[7],A41x_c[7],A41x_c[7],A41x_c[7],A41x_c}*{W41x[7],W41x[7],W41x[7],W41x[7],W41x[7],W41x[7],W41x[7],W41x[7],W41x};
	assign sum42x = {A42x_c[7],A42x_c[7],A42x_c[7],A42x_c[7],A42x_c[7],A42x_c[7],A42x_c[7],A42x_c[7],A42x_c}*{W42x[7],W42x[7],W42x[7],W42x[7],W42x[7],W42x[7],W42x[7],W42x[7],W42x};
	assign sum43x = {A43x_c[7],A43x_c[7],A43x_c[7],A43x_c[7],A43x_c[7],A43x_c[7],A43x_c[7],A43x_c[7],A43x_c}*{W43x[7],W43x[7],W43x[7],W43x[7],W43x[7],W43x[7],W43x[7],W43x[7],W43x};
	assign sum44x = {A44x_c[7],A44x_c[7],A44x_c[7],A44x_c[7],A44x_c[7],A44x_c[7],A44x_c[7],A44x_c[7],A44x_c}*{W44x[7],W44x[7],W44x[7],W44x[7],W44x[7],W44x[7],W44x[7],W44x[7],W44x};
	assign sum45x = {A45x_c[7],A45x_c[7],A45x_c[7],A45x_c[7],A45x_c[7],A45x_c[7],A45x_c[7],A45x_c[7],A45x_c}*{W45x[7],W45x[7],W45x[7],W45x[7],W45x[7],W45x[7],W45x[7],W45x[7],W45x};
	assign sum46x = {A46x_c[7],A46x_c[7],A46x_c[7],A46x_c[7],A46x_c[7],A46x_c[7],A46x_c[7],A46x_c[7],A46x_c}*{W46x[7],W46x[7],W46x[7],W46x[7],W46x[7],W46x[7],W46x[7],W46x[7],W46x};
	assign sum47x = {A47x_c[7],A47x_c[7],A47x_c[7],A47x_c[7],A47x_c[7],A47x_c[7],A47x_c[7],A47x_c[7],A47x_c}*{W47x[7],W47x[7],W47x[7],W47x[7],W47x[7],W47x[7],W47x[7],W47x[7],W47x};
	assign sum48x = {A48x_c[7],A48x_c[7],A48x_c[7],A48x_c[7],A48x_c[7],A48x_c[7],A48x_c[7],A48x_c[7],A48x_c}*{W48x[7],W48x[7],W48x[7],W48x[7],W48x[7],W48x[7],W48x[7],W48x[7],W48x};
	assign sum49x = {A49x_c[7],A49x_c[7],A49x_c[7],A49x_c[7],A49x_c[7],A49x_c[7],A49x_c[7],A49x_c[7],A49x_c}*{W49x[7],W49x[7],W49x[7],W49x[7],W49x[7],W49x[7],W49x[7],W49x[7],W49x};
	assign sum50x = {A50x_c[7],A50x_c[7],A50x_c[7],A50x_c[7],A50x_c[7],A50x_c[7],A50x_c[7],A50x_c[7],A50x_c}*{W50x[7],W50x[7],W50x[7],W50x[7],W50x[7],W50x[7],W50x[7],W50x[7],W50x};
	assign sum51x = {A51x_c[7],A51x_c[7],A51x_c[7],A51x_c[7],A51x_c[7],A51x_c[7],A51x_c[7],A51x_c[7],A51x_c}*{W51x[7],W51x[7],W51x[7],W51x[7],W51x[7],W51x[7],W51x[7],W51x[7],W51x};
	assign sum52x = {A52x_c[7],A52x_c[7],A52x_c[7],A52x_c[7],A52x_c[7],A52x_c[7],A52x_c[7],A52x_c[7],A52x_c}*{W52x[7],W52x[7],W52x[7],W52x[7],W52x[7],W52x[7],W52x[7],W52x[7],W52x};
	assign sum53x = {A53x_c[7],A53x_c[7],A53x_c[7],A53x_c[7],A53x_c[7],A53x_c[7],A53x_c[7],A53x_c[7],A53x_c}*{W53x[7],W53x[7],W53x[7],W53x[7],W53x[7],W53x[7],W53x[7],W53x[7],W53x};
	assign sum54x = {A54x_c[7],A54x_c[7],A54x_c[7],A54x_c[7],A54x_c[7],A54x_c[7],A54x_c[7],A54x_c[7],A54x_c}*{W54x[7],W54x[7],W54x[7],W54x[7],W54x[7],W54x[7],W54x[7],W54x[7],W54x};
	assign sum55x = {A55x_c[7],A55x_c[7],A55x_c[7],A55x_c[7],A55x_c[7],A55x_c[7],A55x_c[7],A55x_c[7],A55x_c}*{W55x[7],W55x[7],W55x[7],W55x[7],W55x[7],W55x[7],W55x[7],W55x[7],W55x};
	assign sum56x = {A56x_c[7],A56x_c[7],A56x_c[7],A56x_c[7],A56x_c[7],A56x_c[7],A56x_c[7],A56x_c[7],A56x_c}*{W56x[7],W56x[7],W56x[7],W56x[7],W56x[7],W56x[7],W56x[7],W56x[7],W56x};
	assign sum57x = {A57x_c[7],A57x_c[7],A57x_c[7],A57x_c[7],A57x_c[7],A57x_c[7],A57x_c[7],A57x_c[7],A57x_c}*{W57x[7],W57x[7],W57x[7],W57x[7],W57x[7],W57x[7],W57x[7],W57x[7],W57x};
	assign sum58x = {A58x_c[7],A58x_c[7],A58x_c[7],A58x_c[7],A58x_c[7],A58x_c[7],A58x_c[7],A58x_c[7],A58x_c}*{W58x[7],W58x[7],W58x[7],W58x[7],W58x[7],W58x[7],W58x[7],W58x[7],W58x};
	assign sum59x = {A59x_c[7],A59x_c[7],A59x_c[7],A59x_c[7],A59x_c[7],A59x_c[7],A59x_c[7],A59x_c[7],A59x_c}*{W59x[7],W59x[7],W59x[7],W59x[7],W59x[7],W59x[7],W59x[7],W59x[7],W59x};
	assign sum60x = {A60x_c[7],A60x_c[7],A60x_c[7],A60x_c[7],A60x_c[7],A60x_c[7],A60x_c[7],A60x_c[7],A60x_c}*{W60x[7],W60x[7],W60x[7],W60x[7],W60x[7],W60x[7],W60x[7],W60x[7],W60x};
	assign sum61x = {A61x_c[7],A61x_c[7],A61x_c[7],A61x_c[7],A61x_c[7],A61x_c[7],A61x_c[7],A61x_c[7],A61x_c}*{W61x[7],W61x[7],W61x[7],W61x[7],W61x[7],W61x[7],W61x[7],W61x[7],W61x};
	assign sum62x = {A62x_c[7],A62x_c[7],A62x_c[7],A62x_c[7],A62x_c[7],A62x_c[7],A62x_c[7],A62x_c[7],A62x_c}*{W62x[7],W62x[7],W62x[7],W62x[7],W62x[7],W62x[7],W62x[7],W62x[7],W62x};
	assign sum63x = {A63x_c[7],A63x_c[7],A63x_c[7],A63x_c[7],A63x_c[7],A63x_c[7],A63x_c[7],A63x_c[7],A63x_c}*{W63x[7],W63x[7],W63x[7],W63x[7],W63x[7],W63x[7],W63x[7],W63x[7],W63x};
	assign sum64x = {A64x_c[7],A64x_c[7],A64x_c[7],A64x_c[7],A64x_c[7],A64x_c[7],A64x_c[7],A64x_c[7],A64x_c}*{W64x[7],W64x[7],W64x[7],W64x[7],W64x[7],W64x[7],W64x[7],W64x[7],W64x};
	assign sum65x = {A65x_c[7],A65x_c[7],A65x_c[7],A65x_c[7],A65x_c[7],A65x_c[7],A65x_c[7],A65x_c[7],A65x_c}*{W65x[7],W65x[7],W65x[7],W65x[7],W65x[7],W65x[7],W65x[7],W65x[7],W65x};
	assign sum66x = {A66x_c[7],A66x_c[7],A66x_c[7],A66x_c[7],A66x_c[7],A66x_c[7],A66x_c[7],A66x_c[7],A66x_c}*{W66x[7],W66x[7],W66x[7],W66x[7],W66x[7],W66x[7],W66x[7],W66x[7],W66x};
	assign sum67x = {A67x_c[7],A67x_c[7],A67x_c[7],A67x_c[7],A67x_c[7],A67x_c[7],A67x_c[7],A67x_c[7],A67x_c}*{W67x[7],W67x[7],W67x[7],W67x[7],W67x[7],W67x[7],W67x[7],W67x[7],W67x};
	assign sum68x = {A68x_c[7],A68x_c[7],A68x_c[7],A68x_c[7],A68x_c[7],A68x_c[7],A68x_c[7],A68x_c[7],A68x_c}*{W68x[7],W68x[7],W68x[7],W68x[7],W68x[7],W68x[7],W68x[7],W68x[7],W68x};
	assign sum69x = {A69x_c[7],A69x_c[7],A69x_c[7],A69x_c[7],A69x_c[7],A69x_c[7],A69x_c[7],A69x_c[7],A69x_c}*{W69x[7],W69x[7],W69x[7],W69x[7],W69x[7],W69x[7],W69x[7],W69x[7],W69x};
	assign sum70x = {A70x_c[7],A70x_c[7],A70x_c[7],A70x_c[7],A70x_c[7],A70x_c[7],A70x_c[7],A70x_c[7],A70x_c}*{W70x[7],W70x[7],W70x[7],W70x[7],W70x[7],W70x[7],W70x[7],W70x[7],W70x};
	assign sum71x = {A71x_c[7],A71x_c[7],A71x_c[7],A71x_c[7],A71x_c[7],A71x_c[7],A71x_c[7],A71x_c[7],A71x_c}*{W71x[7],W71x[7],W71x[7],W71x[7],W71x[7],W71x[7],W71x[7],W71x[7],W71x};
	assign sum72x = {A72x_c[7],A72x_c[7],A72x_c[7],A72x_c[7],A72x_c[7],A72x_c[7],A72x_c[7],A72x_c[7],A72x_c}*{W72x[7],W72x[7],W72x[7],W72x[7],W72x[7],W72x[7],W72x[7],W72x[7],W72x};
	assign sum73x = {A73x_c[7],A73x_c[7],A73x_c[7],A73x_c[7],A73x_c[7],A73x_c[7],A73x_c[7],A73x_c[7],A73x_c}*{W73x[7],W73x[7],W73x[7],W73x[7],W73x[7],W73x[7],W73x[7],W73x[7],W73x};
	assign sum74x = {A74x_c[7],A74x_c[7],A74x_c[7],A74x_c[7],A74x_c[7],A74x_c[7],A74x_c[7],A74x_c[7],A74x_c}*{W74x[7],W74x[7],W74x[7],W74x[7],W74x[7],W74x[7],W74x[7],W74x[7],W74x};
	assign sum75x = {A75x_c[7],A75x_c[7],A75x_c[7],A75x_c[7],A75x_c[7],A75x_c[7],A75x_c[7],A75x_c[7],A75x_c}*{W75x[7],W75x[7],W75x[7],W75x[7],W75x[7],W75x[7],W75x[7],W75x[7],W75x};
	assign sum76x = {A76x_c[7],A76x_c[7],A76x_c[7],A76x_c[7],A76x_c[7],A76x_c[7],A76x_c[7],A76x_c[7],A76x_c}*{W76x[7],W76x[7],W76x[7],W76x[7],W76x[7],W76x[7],W76x[7],W76x[7],W76x};
	assign sum77x = {A77x_c[7],A77x_c[7],A77x_c[7],A77x_c[7],A77x_c[7],A77x_c[7],A77x_c[7],A77x_c[7],A77x_c}*{W77x[7],W77x[7],W77x[7],W77x[7],W77x[7],W77x[7],W77x[7],W77x[7],W77x};
	assign sum78x = {A78x_c[7],A78x_c[7],A78x_c[7],A78x_c[7],A78x_c[7],A78x_c[7],A78x_c[7],A78x_c[7],A78x_c}*{W78x[7],W78x[7],W78x[7],W78x[7],W78x[7],W78x[7],W78x[7],W78x[7],W78x};
	assign sum79x = {A79x_c[7],A79x_c[7],A79x_c[7],A79x_c[7],A79x_c[7],A79x_c[7],A79x_c[7],A79x_c[7],A79x_c}*{W79x[7],W79x[7],W79x[7],W79x[7],W79x[7],W79x[7],W79x[7],W79x[7],W79x};
	assign sum80x = {A80x_c[7],A80x_c[7],A80x_c[7],A80x_c[7],A80x_c[7],A80x_c[7],A80x_c[7],A80x_c[7],A80x_c}*{W80x[7],W80x[7],W80x[7],W80x[7],W80x[7],W80x[7],W80x[7],W80x[7],W80x};
	assign sum81x = {A81x_c[7],A81x_c[7],A81x_c[7],A81x_c[7],A81x_c[7],A81x_c[7],A81x_c[7],A81x_c[7],A81x_c}*{W81x[7],W81x[7],W81x[7],W81x[7],W81x[7],W81x[7],W81x[7],W81x[7],W81x};
	assign sum82x = {A82x_c[7],A82x_c[7],A82x_c[7],A82x_c[7],A82x_c[7],A82x_c[7],A82x_c[7],A82x_c[7],A82x_c}*{W82x[7],W82x[7],W82x[7],W82x[7],W82x[7],W82x[7],W82x[7],W82x[7],W82x};
	assign sum83x = {A83x_c[7],A83x_c[7],A83x_c[7],A83x_c[7],A83x_c[7],A83x_c[7],A83x_c[7],A83x_c[7],A83x_c}*{W83x[7],W83x[7],W83x[7],W83x[7],W83x[7],W83x[7],W83x[7],W83x[7],W83x};
	assign sum84x = {A84x_c[7],A84x_c[7],A84x_c[7],A84x_c[7],A84x_c[7],A84x_c[7],A84x_c[7],A84x_c[7],A84x_c}*{W84x[7],W84x[7],W84x[7],W84x[7],W84x[7],W84x[7],W84x[7],W84x[7],W84x};
	assign sum85x = {A85x_c[7],A85x_c[7],A85x_c[7],A85x_c[7],A85x_c[7],A85x_c[7],A85x_c[7],A85x_c[7],A85x_c}*{W85x[7],W85x[7],W85x[7],W85x[7],W85x[7],W85x[7],W85x[7],W85x[7],W85x};
	assign sum86x = {A86x_c[7],A86x_c[7],A86x_c[7],A86x_c[7],A86x_c[7],A86x_c[7],A86x_c[7],A86x_c[7],A86x_c}*{W86x[7],W86x[7],W86x[7],W86x[7],W86x[7],W86x[7],W86x[7],W86x[7],W86x};
	assign sum87x = {A87x_c[7],A87x_c[7],A87x_c[7],A87x_c[7],A87x_c[7],A87x_c[7],A87x_c[7],A87x_c[7],A87x_c}*{W87x[7],W87x[7],W87x[7],W87x[7],W87x[7],W87x[7],W87x[7],W87x[7],W87x};
	assign sum88x = {A88x_c[7],A88x_c[7],A88x_c[7],A88x_c[7],A88x_c[7],A88x_c[7],A88x_c[7],A88x_c[7],A88x_c}*{W88x[7],W88x[7],W88x[7],W88x[7],W88x[7],W88x[7],W88x[7],W88x[7],W88x};
	assign sum89x = {A89x_c[7],A89x_c[7],A89x_c[7],A89x_c[7],A89x_c[7],A89x_c[7],A89x_c[7],A89x_c[7],A89x_c}*{W89x[7],W89x[7],W89x[7],W89x[7],W89x[7],W89x[7],W89x[7],W89x[7],W89x};
	assign sum90x = {A90x_c[7],A90x_c[7],A90x_c[7],A90x_c[7],A90x_c[7],A90x_c[7],A90x_c[7],A90x_c[7],A90x_c}*{W90x[7],W90x[7],W90x[7],W90x[7],W90x[7],W90x[7],W90x[7],W90x[7],W90x};
	assign sum91x = {A91x_c[7],A91x_c[7],A91x_c[7],A91x_c[7],A91x_c[7],A91x_c[7],A91x_c[7],A91x_c[7],A91x_c}*{W91x[7],W91x[7],W91x[7],W91x[7],W91x[7],W91x[7],W91x[7],W91x[7],W91x};
	assign sum92x = {A92x_c[7],A92x_c[7],A92x_c[7],A92x_c[7],A92x_c[7],A92x_c[7],A92x_c[7],A92x_c[7],A92x_c}*{W92x[7],W92x[7],W92x[7],W92x[7],W92x[7],W92x[7],W92x[7],W92x[7],W92x};
	assign sum93x = {A93x_c[7],A93x_c[7],A93x_c[7],A93x_c[7],A93x_c[7],A93x_c[7],A93x_c[7],A93x_c[7],A93x_c}*{W93x[7],W93x[7],W93x[7],W93x[7],W93x[7],W93x[7],W93x[7],W93x[7],W93x};
	assign sum94x = {A94x_c[7],A94x_c[7],A94x_c[7],A94x_c[7],A94x_c[7],A94x_c[7],A94x_c[7],A94x_c[7],A94x_c}*{W94x[7],W94x[7],W94x[7],W94x[7],W94x[7],W94x[7],W94x[7],W94x[7],W94x};
	assign sum95x = {A95x_c[7],A95x_c[7],A95x_c[7],A95x_c[7],A95x_c[7],A95x_c[7],A95x_c[7],A95x_c[7],A95x_c}*{W95x[7],W95x[7],W95x[7],W95x[7],W95x[7],W95x[7],W95x[7],W95x[7],W95x};
	assign sum96x = {A96x_c[7],A96x_c[7],A96x_c[7],A96x_c[7],A96x_c[7],A96x_c[7],A96x_c[7],A96x_c[7],A96x_c}*{W96x[7],W96x[7],W96x[7],W96x[7],W96x[7],W96x[7],W96x[7],W96x[7],W96x};
	assign sum97x = {A97x_c[7],A97x_c[7],A97x_c[7],A97x_c[7],A97x_c[7],A97x_c[7],A97x_c[7],A97x_c[7],A97x_c}*{W97x[7],W97x[7],W97x[7],W97x[7],W97x[7],W97x[7],W97x[7],W97x[7],W97x};
	assign sum98x = {A98x_c[7],A98x_c[7],A98x_c[7],A98x_c[7],A98x_c[7],A98x_c[7],A98x_c[7],A98x_c[7],A98x_c}*{W98x[7],W98x[7],W98x[7],W98x[7],W98x[7],W98x[7],W98x[7],W98x[7],W98x};
	assign sum99x = {A99x_c[7],A99x_c[7],A99x_c[7],A99x_c[7],A99x_c[7],A99x_c[7],A99x_c[7],A99x_c[7],A99x_c}*{W99x[7],W99x[7],W99x[7],W99x[7],W99x[7],W99x[7],W99x[7],W99x[7],W99x};
	assign sum100x = {A100x_c[7],A100x_c[7],A100x_c[7],A100x_c[7],A100x_c[7],A100x_c[7],A100x_c[7],A100x_c[7],A100x_c}*{W100x[7],W100x[7],W100x[7],W100x[7],W100x[7],W100x[7],W100x[7],W100x[7],W100x};
	assign sum101x = {A101x_c[7],A101x_c[7],A101x_c[7],A101x_c[7],A101x_c[7],A101x_c[7],A101x_c[7],A101x_c[7],A101x_c}*{W101x[7],W101x[7],W101x[7],W101x[7],W101x[7],W101x[7],W101x[7],W101x[7],W101x};
	assign sum102x = {A102x_c[7],A102x_c[7],A102x_c[7],A102x_c[7],A102x_c[7],A102x_c[7],A102x_c[7],A102x_c[7],A102x_c}*{W102x[7],W102x[7],W102x[7],W102x[7],W102x[7],W102x[7],W102x[7],W102x[7],W102x};
	assign sum103x = {A103x_c[7],A103x_c[7],A103x_c[7],A103x_c[7],A103x_c[7],A103x_c[7],A103x_c[7],A103x_c[7],A103x_c}*{W103x[7],W103x[7],W103x[7],W103x[7],W103x[7],W103x[7],W103x[7],W103x[7],W103x};
	assign sum104x = {A104x_c[7],A104x_c[7],A104x_c[7],A104x_c[7],A104x_c[7],A104x_c[7],A104x_c[7],A104x_c[7],A104x_c}*{W104x[7],W104x[7],W104x[7],W104x[7],W104x[7],W104x[7],W104x[7],W104x[7],W104x};
	assign sum105x = {A105x_c[7],A105x_c[7],A105x_c[7],A105x_c[7],A105x_c[7],A105x_c[7],A105x_c[7],A105x_c[7],A105x_c}*{W105x[7],W105x[7],W105x[7],W105x[7],W105x[7],W105x[7],W105x[7],W105x[7],W105x};
	assign sum106x = {A106x_c[7],A106x_c[7],A106x_c[7],A106x_c[7],A106x_c[7],A106x_c[7],A106x_c[7],A106x_c[7],A106x_c}*{W106x[7],W106x[7],W106x[7],W106x[7],W106x[7],W106x[7],W106x[7],W106x[7],W106x};
	assign sum107x = {A107x_c[7],A107x_c[7],A107x_c[7],A107x_c[7],A107x_c[7],A107x_c[7],A107x_c[7],A107x_c[7],A107x_c}*{W107x[7],W107x[7],W107x[7],W107x[7],W107x[7],W107x[7],W107x[7],W107x[7],W107x};
	assign sum108x = {A108x_c[7],A108x_c[7],A108x_c[7],A108x_c[7],A108x_c[7],A108x_c[7],A108x_c[7],A108x_c[7],A108x_c}*{W108x[7],W108x[7],W108x[7],W108x[7],W108x[7],W108x[7],W108x[7],W108x[7],W108x};
	assign sum109x = {A109x_c[7],A109x_c[7],A109x_c[7],A109x_c[7],A109x_c[7],A109x_c[7],A109x_c[7],A109x_c[7],A109x_c}*{W109x[7],W109x[7],W109x[7],W109x[7],W109x[7],W109x[7],W109x[7],W109x[7],W109x};
	assign sum110x = {A110x_c[7],A110x_c[7],A110x_c[7],A110x_c[7],A110x_c[7],A110x_c[7],A110x_c[7],A110x_c[7],A110x_c}*{W110x[7],W110x[7],W110x[7],W110x[7],W110x[7],W110x[7],W110x[7],W110x[7],W110x};
	assign sum111x = {A111x_c[7],A111x_c[7],A111x_c[7],A111x_c[7],A111x_c[7],A111x_c[7],A111x_c[7],A111x_c[7],A111x_c}*{W111x[7],W111x[7],W111x[7],W111x[7],W111x[7],W111x[7],W111x[7],W111x[7],W111x};
	assign sum112x = {A112x_c[7],A112x_c[7],A112x_c[7],A112x_c[7],A112x_c[7],A112x_c[7],A112x_c[7],A112x_c[7],A112x_c}*{W112x[7],W112x[7],W112x[7],W112x[7],W112x[7],W112x[7],W112x[7],W112x[7],W112x};
	assign sum113x = {A113x_c[7],A113x_c[7],A113x_c[7],A113x_c[7],A113x_c[7],A113x_c[7],A113x_c[7],A113x_c[7],A113x_c}*{W113x[7],W113x[7],W113x[7],W113x[7],W113x[7],W113x[7],W113x[7],W113x[7],W113x};
	assign sum114x = {A114x_c[7],A114x_c[7],A114x_c[7],A114x_c[7],A114x_c[7],A114x_c[7],A114x_c[7],A114x_c[7],A114x_c}*{W114x[7],W114x[7],W114x[7],W114x[7],W114x[7],W114x[7],W114x[7],W114x[7],W114x};
	assign sum115x = {A115x_c[7],A115x_c[7],A115x_c[7],A115x_c[7],A115x_c[7],A115x_c[7],A115x_c[7],A115x_c[7],A115x_c}*{W115x[7],W115x[7],W115x[7],W115x[7],W115x[7],W115x[7],W115x[7],W115x[7],W115x};
	assign sum116x = {A116x_c[7],A116x_c[7],A116x_c[7],A116x_c[7],A116x_c[7],A116x_c[7],A116x_c[7],A116x_c[7],A116x_c}*{W116x[7],W116x[7],W116x[7],W116x[7],W116x[7],W116x[7],W116x[7],W116x[7],W116x};
	assign sum117x = {A117x_c[7],A117x_c[7],A117x_c[7],A117x_c[7],A117x_c[7],A117x_c[7],A117x_c[7],A117x_c[7],A117x_c}*{W117x[7],W117x[7],W117x[7],W117x[7],W117x[7],W117x[7],W117x[7],W117x[7],W117x};
	assign sum118x = {A118x_c[7],A118x_c[7],A118x_c[7],A118x_c[7],A118x_c[7],A118x_c[7],A118x_c[7],A118x_c[7],A118x_c}*{W118x[7],W118x[7],W118x[7],W118x[7],W118x[7],W118x[7],W118x[7],W118x[7],W118x};
	assign sum119x = {A119x_c[7],A119x_c[7],A119x_c[7],A119x_c[7],A119x_c[7],A119x_c[7],A119x_c[7],A119x_c[7],A119x_c}*{W119x[7],W119x[7],W119x[7],W119x[7],W119x[7],W119x[7],W119x[7],W119x[7],W119x};
	assign sum120x = {A120x_c[7],A120x_c[7],A120x_c[7],A120x_c[7],A120x_c[7],A120x_c[7],A120x_c[7],A120x_c[7],A120x_c}*{W120x[7],W120x[7],W120x[7],W120x[7],W120x[7],W120x[7],W120x[7],W120x[7],W120x};
	assign sum121x = {A121x_c[7],A121x_c[7],A121x_c[7],A121x_c[7],A121x_c[7],A121x_c[7],A121x_c[7],A121x_c[7],A121x_c}*{W121x[7],W121x[7],W121x[7],W121x[7],W121x[7],W121x[7],W121x[7],W121x[7],W121x};
	assign sum122x = {A122x_c[7],A122x_c[7],A122x_c[7],A122x_c[7],A122x_c[7],A122x_c[7],A122x_c[7],A122x_c[7],A122x_c}*{W122x[7],W122x[7],W122x[7],W122x[7],W122x[7],W122x[7],W122x[7],W122x[7],W122x};
	assign sum123x = {A123x_c[7],A123x_c[7],A123x_c[7],A123x_c[7],A123x_c[7],A123x_c[7],A123x_c[7],A123x_c[7],A123x_c}*{W123x[7],W123x[7],W123x[7],W123x[7],W123x[7],W123x[7],W123x[7],W123x[7],W123x};
	assign sum124x = {A124x_c[7],A124x_c[7],A124x_c[7],A124x_c[7],A124x_c[7],A124x_c[7],A124x_c[7],A124x_c[7],A124x_c}*{W124x[7],W124x[7],W124x[7],W124x[7],W124x[7],W124x[7],W124x[7],W124x[7],W124x};
	assign sum125x = {A125x_c[7],A125x_c[7],A125x_c[7],A125x_c[7],A125x_c[7],A125x_c[7],A125x_c[7],A125x_c[7],A125x_c}*{W125x[7],W125x[7],W125x[7],W125x[7],W125x[7],W125x[7],W125x[7],W125x[7],W125x};
	assign sum126x = {A126x_c[7],A126x_c[7],A126x_c[7],A126x_c[7],A126x_c[7],A126x_c[7],A126x_c[7],A126x_c[7],A126x_c}*{W126x[7],W126x[7],W126x[7],W126x[7],W126x[7],W126x[7],W126x[7],W126x[7],W126x};
	assign sum127x = {A127x_c[7],A127x_c[7],A127x_c[7],A127x_c[7],A127x_c[7],A127x_c[7],A127x_c[7],A127x_c[7],A127x_c}*{W127x[7],W127x[7],W127x[7],W127x[7],W127x[7],W127x[7],W127x[7],W127x[7],W127x};
	assign sum128x = {A128x_c[7],A128x_c[7],A128x_c[7],A128x_c[7],A128x_c[7],A128x_c[7],A128x_c[7],A128x_c[7],A128x_c}*{W128x[7],W128x[7],W128x[7],W128x[7],W128x[7],W128x[7],W128x[7],W128x[7],W128x};
	assign sum129x = {A129x_c[7],A129x_c[7],A129x_c[7],A129x_c[7],A129x_c[7],A129x_c[7],A129x_c[7],A129x_c[7],A129x_c}*{W129x[7],W129x[7],W129x[7],W129x[7],W129x[7],W129x[7],W129x[7],W129x[7],W129x};
	assign sum130x = {A130x_c[7],A130x_c[7],A130x_c[7],A130x_c[7],A130x_c[7],A130x_c[7],A130x_c[7],A130x_c[7],A130x_c}*{W130x[7],W130x[7],W130x[7],W130x[7],W130x[7],W130x[7],W130x[7],W130x[7],W130x};
	assign sum131x = {A131x_c[7],A131x_c[7],A131x_c[7],A131x_c[7],A131x_c[7],A131x_c[7],A131x_c[7],A131x_c[7],A131x_c}*{W131x[7],W131x[7],W131x[7],W131x[7],W131x[7],W131x[7],W131x[7],W131x[7],W131x};
	assign sum132x = {A132x_c[7],A132x_c[7],A132x_c[7],A132x_c[7],A132x_c[7],A132x_c[7],A132x_c[7],A132x_c[7],A132x_c}*{W132x[7],W132x[7],W132x[7],W132x[7],W132x[7],W132x[7],W132x[7],W132x[7],W132x};
	assign sum133x = {A133x_c[7],A133x_c[7],A133x_c[7],A133x_c[7],A133x_c[7],A133x_c[7],A133x_c[7],A133x_c[7],A133x_c}*{W133x[7],W133x[7],W133x[7],W133x[7],W133x[7],W133x[7],W133x[7],W133x[7],W133x};
	assign sum134x = {A134x_c[7],A134x_c[7],A134x_c[7],A134x_c[7],A134x_c[7],A134x_c[7],A134x_c[7],A134x_c[7],A134x_c}*{W134x[7],W134x[7],W134x[7],W134x[7],W134x[7],W134x[7],W134x[7],W134x[7],W134x};
	assign sum135x = {A135x_c[7],A135x_c[7],A135x_c[7],A135x_c[7],A135x_c[7],A135x_c[7],A135x_c[7],A135x_c[7],A135x_c}*{W135x[7],W135x[7],W135x[7],W135x[7],W135x[7],W135x[7],W135x[7],W135x[7],W135x};
	assign sum136x = {A136x_c[7],A136x_c[7],A136x_c[7],A136x_c[7],A136x_c[7],A136x_c[7],A136x_c[7],A136x_c[7],A136x_c}*{W136x[7],W136x[7],W136x[7],W136x[7],W136x[7],W136x[7],W136x[7],W136x[7],W136x};
	assign sum137x = {A137x_c[7],A137x_c[7],A137x_c[7],A137x_c[7],A137x_c[7],A137x_c[7],A137x_c[7],A137x_c[7],A137x_c}*{W137x[7],W137x[7],W137x[7],W137x[7],W137x[7],W137x[7],W137x[7],W137x[7],W137x};
	assign sum138x = {A138x_c[7],A138x_c[7],A138x_c[7],A138x_c[7],A138x_c[7],A138x_c[7],A138x_c[7],A138x_c[7],A138x_c}*{W138x[7],W138x[7],W138x[7],W138x[7],W138x[7],W138x[7],W138x[7],W138x[7],W138x};
	assign sum139x = {A139x_c[7],A139x_c[7],A139x_c[7],A139x_c[7],A139x_c[7],A139x_c[7],A139x_c[7],A139x_c[7],A139x_c}*{W139x[7],W139x[7],W139x[7],W139x[7],W139x[7],W139x[7],W139x[7],W139x[7],W139x};
	assign sum140x = {A140x_c[7],A140x_c[7],A140x_c[7],A140x_c[7],A140x_c[7],A140x_c[7],A140x_c[7],A140x_c[7],A140x_c}*{W140x[7],W140x[7],W140x[7],W140x[7],W140x[7],W140x[7],W140x[7],W140x[7],W140x};
	assign sum141x = {A141x_c[7],A141x_c[7],A141x_c[7],A141x_c[7],A141x_c[7],A141x_c[7],A141x_c[7],A141x_c[7],A141x_c}*{W141x[7],W141x[7],W141x[7],W141x[7],W141x[7],W141x[7],W141x[7],W141x[7],W141x};
	assign sum142x = {A142x_c[7],A142x_c[7],A142x_c[7],A142x_c[7],A142x_c[7],A142x_c[7],A142x_c[7],A142x_c[7],A142x_c}*{W142x[7],W142x[7],W142x[7],W142x[7],W142x[7],W142x[7],W142x[7],W142x[7],W142x};
	assign sum143x = {A143x_c[7],A143x_c[7],A143x_c[7],A143x_c[7],A143x_c[7],A143x_c[7],A143x_c[7],A143x_c[7],A143x_c}*{W143x[7],W143x[7],W143x[7],W143x[7],W143x[7],W143x[7],W143x[7],W143x[7],W143x};
	assign sum144x = {A144x_c[7],A144x_c[7],A144x_c[7],A144x_c[7],A144x_c[7],A144x_c[7],A144x_c[7],A144x_c[7],A144x_c}*{W144x[7],W144x[7],W144x[7],W144x[7],W144x[7],W144x[7],W144x[7],W144x[7],W144x};
	assign sum145x = {A145x_c[7],A145x_c[7],A145x_c[7],A145x_c[7],A145x_c[7],A145x_c[7],A145x_c[7],A145x_c[7],A145x_c}*{W145x[7],W145x[7],W145x[7],W145x[7],W145x[7],W145x[7],W145x[7],W145x[7],W145x};
	assign sum146x = {A146x_c[7],A146x_c[7],A146x_c[7],A146x_c[7],A146x_c[7],A146x_c[7],A146x_c[7],A146x_c[7],A146x_c}*{W146x[7],W146x[7],W146x[7],W146x[7],W146x[7],W146x[7],W146x[7],W146x[7],W146x};
	assign sum147x = {A147x_c[7],A147x_c[7],A147x_c[7],A147x_c[7],A147x_c[7],A147x_c[7],A147x_c[7],A147x_c[7],A147x_c}*{W147x[7],W147x[7],W147x[7],W147x[7],W147x[7],W147x[7],W147x[7],W147x[7],W147x};
	assign sum148x = {A148x_c[7],A148x_c[7],A148x_c[7],A148x_c[7],A148x_c[7],A148x_c[7],A148x_c[7],A148x_c[7],A148x_c}*{W148x[7],W148x[7],W148x[7],W148x[7],W148x[7],W148x[7],W148x[7],W148x[7],W148x};
	assign sum149x = {A149x_c[7],A149x_c[7],A149x_c[7],A149x_c[7],A149x_c[7],A149x_c[7],A149x_c[7],A149x_c[7],A149x_c}*{W149x[7],W149x[7],W149x[7],W149x[7],W149x[7],W149x[7],W149x[7],W149x[7],W149x};
	assign sum150x = {A150x_c[7],A150x_c[7],A150x_c[7],A150x_c[7],A150x_c[7],A150x_c[7],A150x_c[7],A150x_c[7],A150x_c}*{W150x[7],W150x[7],W150x[7],W150x[7],W150x[7],W150x[7],W150x[7],W150x[7],W150x};
	assign sum151x = {A151x_c[7],A151x_c[7],A151x_c[7],A151x_c[7],A151x_c[7],A151x_c[7],A151x_c[7],A151x_c[7],A151x_c}*{W151x[7],W151x[7],W151x[7],W151x[7],W151x[7],W151x[7],W151x[7],W151x[7],W151x};
	assign sum152x = {A152x_c[7],A152x_c[7],A152x_c[7],A152x_c[7],A152x_c[7],A152x_c[7],A152x_c[7],A152x_c[7],A152x_c}*{W152x[7],W152x[7],W152x[7],W152x[7],W152x[7],W152x[7],W152x[7],W152x[7],W152x};
	assign sum153x = {A153x_c[7],A153x_c[7],A153x_c[7],A153x_c[7],A153x_c[7],A153x_c[7],A153x_c[7],A153x_c[7],A153x_c}*{W153x[7],W153x[7],W153x[7],W153x[7],W153x[7],W153x[7],W153x[7],W153x[7],W153x};
	assign sum154x = {A154x_c[7],A154x_c[7],A154x_c[7],A154x_c[7],A154x_c[7],A154x_c[7],A154x_c[7],A154x_c[7],A154x_c}*{W154x[7],W154x[7],W154x[7],W154x[7],W154x[7],W154x[7],W154x[7],W154x[7],W154x};
	assign sum155x = {A155x_c[7],A155x_c[7],A155x_c[7],A155x_c[7],A155x_c[7],A155x_c[7],A155x_c[7],A155x_c[7],A155x_c}*{W155x[7],W155x[7],W155x[7],W155x[7],W155x[7],W155x[7],W155x[7],W155x[7],W155x};
	assign sum156x = {A156x_c[7],A156x_c[7],A156x_c[7],A156x_c[7],A156x_c[7],A156x_c[7],A156x_c[7],A156x_c[7],A156x_c}*{W156x[7],W156x[7],W156x[7],W156x[7],W156x[7],W156x[7],W156x[7],W156x[7],W156x};
	assign sum157x = {A157x_c[7],A157x_c[7],A157x_c[7],A157x_c[7],A157x_c[7],A157x_c[7],A157x_c[7],A157x_c[7],A157x_c}*{W157x[7],W157x[7],W157x[7],W157x[7],W157x[7],W157x[7],W157x[7],W157x[7],W157x};
	assign sum158x = {A158x_c[7],A158x_c[7],A158x_c[7],A158x_c[7],A158x_c[7],A158x_c[7],A158x_c[7],A158x_c[7],A158x_c}*{W158x[7],W158x[7],W158x[7],W158x[7],W158x[7],W158x[7],W158x[7],W158x[7],W158x};
	assign sum159x = {A159x_c[7],A159x_c[7],A159x_c[7],A159x_c[7],A159x_c[7],A159x_c[7],A159x_c[7],A159x_c[7],A159x_c}*{W159x[7],W159x[7],W159x[7],W159x[7],W159x[7],W159x[7],W159x[7],W159x[7],W159x};
	assign sum160x = {A160x_c[7],A160x_c[7],A160x_c[7],A160x_c[7],A160x_c[7],A160x_c[7],A160x_c[7],A160x_c[7],A160x_c}*{W160x[7],W160x[7],W160x[7],W160x[7],W160x[7],W160x[7],W160x[7],W160x[7],W160x};
	assign sum161x = {A161x_c[7],A161x_c[7],A161x_c[7],A161x_c[7],A161x_c[7],A161x_c[7],A161x_c[7],A161x_c[7],A161x_c}*{W161x[7],W161x[7],W161x[7],W161x[7],W161x[7],W161x[7],W161x[7],W161x[7],W161x};
	assign sum162x = {A162x_c[7],A162x_c[7],A162x_c[7],A162x_c[7],A162x_c[7],A162x_c[7],A162x_c[7],A162x_c[7],A162x_c}*{W162x[7],W162x[7],W162x[7],W162x[7],W162x[7],W162x[7],W162x[7],W162x[7],W162x};
	assign sum163x = {A163x_c[7],A163x_c[7],A163x_c[7],A163x_c[7],A163x_c[7],A163x_c[7],A163x_c[7],A163x_c[7],A163x_c}*{W163x[7],W163x[7],W163x[7],W163x[7],W163x[7],W163x[7],W163x[7],W163x[7],W163x};
	assign sum164x = {A164x_c[7],A164x_c[7],A164x_c[7],A164x_c[7],A164x_c[7],A164x_c[7],A164x_c[7],A164x_c[7],A164x_c}*{W164x[7],W164x[7],W164x[7],W164x[7],W164x[7],W164x[7],W164x[7],W164x[7],W164x};
	assign sum165x = {A165x_c[7],A165x_c[7],A165x_c[7],A165x_c[7],A165x_c[7],A165x_c[7],A165x_c[7],A165x_c[7],A165x_c}*{W165x[7],W165x[7],W165x[7],W165x[7],W165x[7],W165x[7],W165x[7],W165x[7],W165x};
	assign sum166x = {A166x_c[7],A166x_c[7],A166x_c[7],A166x_c[7],A166x_c[7],A166x_c[7],A166x_c[7],A166x_c[7],A166x_c}*{W166x[7],W166x[7],W166x[7],W166x[7],W166x[7],W166x[7],W166x[7],W166x[7],W166x};
	assign sum167x = {A167x_c[7],A167x_c[7],A167x_c[7],A167x_c[7],A167x_c[7],A167x_c[7],A167x_c[7],A167x_c[7],A167x_c}*{W167x[7],W167x[7],W167x[7],W167x[7],W167x[7],W167x[7],W167x[7],W167x[7],W167x};
	assign sum168x = {A168x_c[7],A168x_c[7],A168x_c[7],A168x_c[7],A168x_c[7],A168x_c[7],A168x_c[7],A168x_c[7],A168x_c}*{W168x[7],W168x[7],W168x[7],W168x[7],W168x[7],W168x[7],W168x[7],W168x[7],W168x};
	assign sum169x = {A169x_c[7],A169x_c[7],A169x_c[7],A169x_c[7],A169x_c[7],A169x_c[7],A169x_c[7],A169x_c[7],A169x_c}*{W169x[7],W169x[7],W169x[7],W169x[7],W169x[7],W169x[7],W169x[7],W169x[7],W169x};
	assign sum170x = {A170x_c[7],A170x_c[7],A170x_c[7],A170x_c[7],A170x_c[7],A170x_c[7],A170x_c[7],A170x_c[7],A170x_c}*{W170x[7],W170x[7],W170x[7],W170x[7],W170x[7],W170x[7],W170x[7],W170x[7],W170x};
	assign sum171x = {A171x_c[7],A171x_c[7],A171x_c[7],A171x_c[7],A171x_c[7],A171x_c[7],A171x_c[7],A171x_c[7],A171x_c}*{W171x[7],W171x[7],W171x[7],W171x[7],W171x[7],W171x[7],W171x[7],W171x[7],W171x};
	assign sum172x = {A172x_c[7],A172x_c[7],A172x_c[7],A172x_c[7],A172x_c[7],A172x_c[7],A172x_c[7],A172x_c[7],A172x_c}*{W172x[7],W172x[7],W172x[7],W172x[7],W172x[7],W172x[7],W172x[7],W172x[7],W172x};
	assign sum173x = {A173x_c[7],A173x_c[7],A173x_c[7],A173x_c[7],A173x_c[7],A173x_c[7],A173x_c[7],A173x_c[7],A173x_c}*{W173x[7],W173x[7],W173x[7],W173x[7],W173x[7],W173x[7],W173x[7],W173x[7],W173x};
	assign sum174x = {A174x_c[7],A174x_c[7],A174x_c[7],A174x_c[7],A174x_c[7],A174x_c[7],A174x_c[7],A174x_c[7],A174x_c}*{W174x[7],W174x[7],W174x[7],W174x[7],W174x[7],W174x[7],W174x[7],W174x[7],W174x};
	assign sum175x = {A175x_c[7],A175x_c[7],A175x_c[7],A175x_c[7],A175x_c[7],A175x_c[7],A175x_c[7],A175x_c[7],A175x_c}*{W175x[7],W175x[7],W175x[7],W175x[7],W175x[7],W175x[7],W175x[7],W175x[7],W175x};
	assign sum176x = {A176x_c[7],A176x_c[7],A176x_c[7],A176x_c[7],A176x_c[7],A176x_c[7],A176x_c[7],A176x_c[7],A176x_c}*{W176x[7],W176x[7],W176x[7],W176x[7],W176x[7],W176x[7],W176x[7],W176x[7],W176x};
	assign sum177x = {A177x_c[7],A177x_c[7],A177x_c[7],A177x_c[7],A177x_c[7],A177x_c[7],A177x_c[7],A177x_c[7],A177x_c}*{W177x[7],W177x[7],W177x[7],W177x[7],W177x[7],W177x[7],W177x[7],W177x[7],W177x};
	assign sum178x = {A178x_c[7],A178x_c[7],A178x_c[7],A178x_c[7],A178x_c[7],A178x_c[7],A178x_c[7],A178x_c[7],A178x_c}*{W178x[7],W178x[7],W178x[7],W178x[7],W178x[7],W178x[7],W178x[7],W178x[7],W178x};
	assign sum179x = {A179x_c[7],A179x_c[7],A179x_c[7],A179x_c[7],A179x_c[7],A179x_c[7],A179x_c[7],A179x_c[7],A179x_c}*{W179x[7],W179x[7],W179x[7],W179x[7],W179x[7],W179x[7],W179x[7],W179x[7],W179x};
	assign sum180x = {A180x_c[7],A180x_c[7],A180x_c[7],A180x_c[7],A180x_c[7],A180x_c[7],A180x_c[7],A180x_c[7],A180x_c}*{W180x[7],W180x[7],W180x[7],W180x[7],W180x[7],W180x[7],W180x[7],W180x[7],W180x};
	assign sum181x = {A181x_c[7],A181x_c[7],A181x_c[7],A181x_c[7],A181x_c[7],A181x_c[7],A181x_c[7],A181x_c[7],A181x_c}*{W181x[7],W181x[7],W181x[7],W181x[7],W181x[7],W181x[7],W181x[7],W181x[7],W181x};
	assign sum182x = {A182x_c[7],A182x_c[7],A182x_c[7],A182x_c[7],A182x_c[7],A182x_c[7],A182x_c[7],A182x_c[7],A182x_c}*{W182x[7],W182x[7],W182x[7],W182x[7],W182x[7],W182x[7],W182x[7],W182x[7],W182x};
	assign sum183x = {A183x_c[7],A183x_c[7],A183x_c[7],A183x_c[7],A183x_c[7],A183x_c[7],A183x_c[7],A183x_c[7],A183x_c}*{W183x[7],W183x[7],W183x[7],W183x[7],W183x[7],W183x[7],W183x[7],W183x[7],W183x};
	assign sum184x = {A184x_c[7],A184x_c[7],A184x_c[7],A184x_c[7],A184x_c[7],A184x_c[7],A184x_c[7],A184x_c[7],A184x_c}*{W184x[7],W184x[7],W184x[7],W184x[7],W184x[7],W184x[7],W184x[7],W184x[7],W184x};
	assign sum185x = {A185x_c[7],A185x_c[7],A185x_c[7],A185x_c[7],A185x_c[7],A185x_c[7],A185x_c[7],A185x_c[7],A185x_c}*{W185x[7],W185x[7],W185x[7],W185x[7],W185x[7],W185x[7],W185x[7],W185x[7],W185x};
	assign sum186x = {A186x_c[7],A186x_c[7],A186x_c[7],A186x_c[7],A186x_c[7],A186x_c[7],A186x_c[7],A186x_c[7],A186x_c}*{W186x[7],W186x[7],W186x[7],W186x[7],W186x[7],W186x[7],W186x[7],W186x[7],W186x};

	always@(posedge clk) begin

		if(reset)
			begin
			N3x<=8'd0;
			sumout<=16'd0;
			A0x_c <= 8'd0;
			A1x_c <= 8'd0;
			A2x_c <= 8'd0;
			A3x_c <= 8'd0;
			A4x_c <= 8'd0;
			A5x_c <= 8'd0;
			A6x_c <= 8'd0;
			A7x_c <= 8'd0;
			A8x_c <= 8'd0;
			A9x_c <= 8'd0;
			A10x_c <= 8'd0;
			A11x_c <= 8'd0;
			A12x_c <= 8'd0;
			A13x_c <= 8'd0;
			A14x_c <= 8'd0;
			A15x_c <= 8'd0;
			A16x_c <= 8'd0;
			A17x_c <= 8'd0;
			A18x_c <= 8'd0;
			A19x_c <= 8'd0;
			A20x_c <= 8'd0;
			A21x_c <= 8'd0;
			A22x_c <= 8'd0;
			A23x_c <= 8'd0;
			A24x_c <= 8'd0;
			A25x_c <= 8'd0;
			A26x_c <= 8'd0;
			A27x_c <= 8'd0;
			A28x_c <= 8'd0;
			A29x_c <= 8'd0;
			A30x_c <= 8'd0;
			A31x_c <= 8'd0;
			A32x_c <= 8'd0;
			A33x_c <= 8'd0;
			A34x_c <= 8'd0;
			A35x_c <= 8'd0;
			A36x_c <= 8'd0;
			A37x_c <= 8'd0;
			A38x_c <= 8'd0;
			A39x_c <= 8'd0;
			A40x_c <= 8'd0;
			A41x_c <= 8'd0;
			A42x_c <= 8'd0;
			A43x_c <= 8'd0;
			A44x_c <= 8'd0;
			A45x_c <= 8'd0;
			A46x_c <= 8'd0;
			A47x_c <= 8'd0;
			A48x_c <= 8'd0;
			A49x_c <= 8'd0;
			A50x_c <= 8'd0;
			A51x_c <= 8'd0;
			A52x_c <= 8'd0;
			A53x_c <= 8'd0;
			A54x_c <= 8'd0;
			A55x_c <= 8'd0;
			A56x_c <= 8'd0;
			A57x_c <= 8'd0;
			A58x_c <= 8'd0;
			A59x_c <= 8'd0;
			A60x_c <= 8'd0;
			A61x_c <= 8'd0;
			A62x_c <= 8'd0;
			A63x_c <= 8'd0;
			A64x_c <= 8'd0;
			A65x_c <= 8'd0;
			A66x_c <= 8'd0;
			A67x_c <= 8'd0;
			A68x_c <= 8'd0;
			A69x_c <= 8'd0;
			A70x_c <= 8'd0;
			A71x_c <= 8'd0;
			A72x_c <= 8'd0;
			A73x_c <= 8'd0;
			A74x_c <= 8'd0;
			A75x_c <= 8'd0;
			A76x_c <= 8'd0;
			A77x_c <= 8'd0;
			A78x_c <= 8'd0;
			A79x_c <= 8'd0;
			A80x_c <= 8'd0;
			A81x_c <= 8'd0;
			A82x_c <= 8'd0;
			A83x_c <= 8'd0;
			A84x_c <= 8'd0;
			A85x_c <= 8'd0;
			A86x_c <= 8'd0;
			A87x_c <= 8'd0;
			A88x_c <= 8'd0;
			A89x_c <= 8'd0;
			A90x_c <= 8'd0;
			A91x_c <= 8'd0;
			A92x_c <= 8'd0;
			A93x_c <= 8'd0;
			A94x_c <= 8'd0;
			A95x_c <= 8'd0;
			A96x_c <= 8'd0;
			A97x_c <= 8'd0;
			A98x_c <= 8'd0;
			A99x_c <= 8'd0;
			A100x_c <= 8'd0;
			A101x_c <= 8'd0;
			A102x_c <= 8'd0;
			A103x_c <= 8'd0;
			A104x_c <= 8'd0;
			A105x_c <= 8'd0;
			A106x_c <= 8'd0;
			A107x_c <= 8'd0;
			A108x_c <= 8'd0;
			A109x_c <= 8'd0;
			A110x_c <= 8'd0;
			A111x_c <= 8'd0;
			A112x_c <= 8'd0;
			A113x_c <= 8'd0;
			A114x_c <= 8'd0;
			A115x_c <= 8'd0;
			A116x_c <= 8'd0;
			A117x_c <= 8'd0;
			A118x_c <= 8'd0;
			A119x_c <= 8'd0;
			A120x_c <= 8'd0;
			A121x_c <= 8'd0;
			A122x_c <= 8'd0;
			A123x_c <= 8'd0;
			A124x_c <= 8'd0;
			A125x_c <= 8'd0;
			A126x_c <= 8'd0;
			A127x_c <= 8'd0;
			A128x_c <= 8'd0;
			A129x_c <= 8'd0;
			A130x_c <= 8'd0;
			A131x_c <= 8'd0;
			A132x_c <= 8'd0;
			A133x_c <= 8'd0;
			A134x_c <= 8'd0;
			A135x_c <= 8'd0;
			A136x_c <= 8'd0;
			A137x_c <= 8'd0;
			A138x_c <= 8'd0;
			A139x_c <= 8'd0;
			A140x_c <= 8'd0;
			A141x_c <= 8'd0;
			A142x_c <= 8'd0;
			A143x_c <= 8'd0;
			A144x_c <= 8'd0;
			A145x_c <= 8'd0;
			A146x_c <= 8'd0;
			A147x_c <= 8'd0;
			A148x_c <= 8'd0;
			A149x_c <= 8'd0;
			A150x_c <= 8'd0;
			A151x_c <= 8'd0;
			A152x_c <= 8'd0;
			A153x_c <= 8'd0;
			A154x_c <= 8'd0;
			A155x_c <= 8'd0;
			A156x_c <= 8'd0;
			A157x_c <= 8'd0;
			A158x_c <= 8'd0;
			A159x_c <= 8'd0;
			A160x_c <= 8'd0;
			A161x_c <= 8'd0;
			A162x_c <= 8'd0;
			A163x_c <= 8'd0;
			A164x_c <= 8'd0;
			A165x_c <= 8'd0;
			A166x_c <= 8'd0;
			A167x_c <= 8'd0;
			A168x_c <= 8'd0;
			A169x_c <= 8'd0;
			A170x_c <= 8'd0;
			A171x_c <= 8'd0;
			A172x_c <= 8'd0;
			A173x_c <= 8'd0;
			A174x_c <= 8'd0;
			A175x_c <= 8'd0;
			A176x_c <= 8'd0;
			A177x_c <= 8'd0;
			A178x_c <= 8'd0;
			A179x_c <= 8'd0;
			A180x_c <= 8'd0;
			A181x_c <= 8'd0;
			A182x_c <= 8'd0;
			A183x_c <= 8'd0;
			A184x_c <= 8'd0;
			A185x_c <= 8'd0;
			A186x_c <= 8'd0;
			end
		else
			begin
			A0x_c <= A0x;
			A1x_c <= A1x;
			A2x_c <= A2x;
			A3x_c <= A3x;
			A4x_c <= A4x;
			A5x_c <= A5x;
			A6x_c <= A6x;
			A7x_c <= A7x;
			A8x_c <= A8x;
			A9x_c <= A9x;
			A10x_c <= A10x;
			A11x_c <= A11x;
			A12x_c <= A12x;
			A13x_c <= A13x;
			A14x_c <= A14x;
			A15x_c <= A15x;
			A16x_c <= A16x;
			A17x_c <= A17x;
			A18x_c <= A18x;
			A19x_c <= A19x;
			A20x_c <= A20x;
			A21x_c <= A21x;
			A22x_c <= A22x;
			A23x_c <= A23x;
			A24x_c <= A24x;
			A25x_c <= A25x;
			A26x_c <= A26x;
			A27x_c <= A27x;
			A28x_c <= A28x;
			A29x_c <= A29x;
			A30x_c <= A30x;
			A31x_c <= A31x;
			A32x_c <= A32x;
			A33x_c <= A33x;
			A34x_c <= A34x;
			A35x_c <= A35x;
			A36x_c <= A36x;
			A37x_c <= A37x;
			A38x_c <= A38x;
			A39x_c <= A39x;
			A40x_c <= A40x;
			A41x_c <= A41x;
			A42x_c <= A42x;
			A43x_c <= A43x;
			A44x_c <= A44x;
			A45x_c <= A45x;
			A46x_c <= A46x;
			A47x_c <= A47x;
			A48x_c <= A48x;
			A49x_c <= A49x;
			A50x_c <= A50x;
			A51x_c <= A51x;
			A52x_c <= A52x;
			A53x_c <= A53x;
			A54x_c <= A54x;
			A55x_c <= A55x;
			A56x_c <= A56x;
			A57x_c <= A57x;
			A58x_c <= A58x;
			A59x_c <= A59x;
			A60x_c <= A60x;
			A61x_c <= A61x;
			A62x_c <= A62x;
			A63x_c <= A63x;
			A64x_c <= A64x;
			A65x_c <= A65x;
			A66x_c <= A66x;
			A67x_c <= A67x;
			A68x_c <= A68x;
			A69x_c <= A69x;
			A70x_c <= A70x;
			A71x_c <= A71x;
			A72x_c <= A72x;
			A73x_c <= A73x;
			A74x_c <= A74x;
			A75x_c <= A75x;
			A76x_c <= A76x;
			A77x_c <= A77x;
			A78x_c <= A78x;
			A79x_c <= A79x;
			A80x_c <= A80x;
			A81x_c <= A81x;
			A82x_c <= A82x;
			A83x_c <= A83x;
			A84x_c <= A84x;
			A85x_c <= A85x;
			A86x_c <= A86x;
			A87x_c <= A87x;
			A88x_c <= A88x;
			A89x_c <= A89x;
			A90x_c <= A90x;
			A91x_c <= A91x;
			A92x_c <= A92x;
			A93x_c <= A93x;
			A94x_c <= A94x;
			A95x_c <= A95x;
			A96x_c <= A96x;
			A97x_c <= A97x;
			A98x_c <= A98x;
			A99x_c <= A99x;
			A100x_c <= A100x;
			A101x_c <= A101x;
			A102x_c <= A102x;
			A103x_c <= A103x;
			A104x_c <= A104x;
			A105x_c <= A105x;
			A106x_c <= A106x;
			A107x_c <= A107x;
			A108x_c <= A108x;
			A109x_c <= A109x;
			A110x_c <= A110x;
			A111x_c <= A111x;
			A112x_c <= A112x;
			A113x_c <= A113x;
			A114x_c <= A114x;
			A115x_c <= A115x;
			A116x_c <= A116x;
			A117x_c <= A117x;
			A118x_c <= A118x;
			A119x_c <= A119x;
			A120x_c <= A120x;
			A121x_c <= A121x;
			A122x_c <= A122x;
			A123x_c <= A123x;
			A124x_c <= A124x;
			A125x_c <= A125x;
			A126x_c <= A126x;
			A127x_c <= A127x;
			A128x_c <= A128x;
			A129x_c <= A129x;
			A130x_c <= A130x;
			A131x_c <= A131x;
			A132x_c <= A132x;
			A133x_c <= A133x;
			A134x_c <= A134x;
			A135x_c <= A135x;
			A136x_c <= A136x;
			A137x_c <= A137x;
			A138x_c <= A138x;
			A139x_c <= A139x;
			A140x_c <= A140x;
			A141x_c <= A141x;
			A142x_c <= A142x;
			A143x_c <= A143x;
			A144x_c <= A144x;
			A145x_c <= A145x;
			A146x_c <= A146x;
			A147x_c <= A147x;
			A148x_c <= A148x;
			A149x_c <= A149x;
			A150x_c <= A150x;
			A151x_c <= A151x;
			A152x_c <= A152x;
			A153x_c <= A153x;
			A154x_c <= A154x;
			A155x_c <= A155x;
			A156x_c <= A156x;
			A157x_c <= A157x;
			A158x_c <= A158x;
			A159x_c <= A159x;
			A160x_c <= A160x;
			A161x_c <= A161x;
			A162x_c <= A162x;
			A163x_c <= A163x;
			A164x_c <= A164x;
			A165x_c <= A165x;
			A166x_c <= A166x;
			A167x_c <= A167x;
			A168x_c <= A168x;
			A169x_c <= A169x;
			A170x_c <= A170x;
			A171x_c <= A171x;
			A172x_c <= A172x;
			A173x_c <= A173x;
			A174x_c <= A174x;
			A175x_c <= A175x;
			A176x_c <= A176x;
			A177x_c <= A177x;
			A178x_c <= A178x;
			A179x_c <= A179x;
			A180x_c <= A180x;
			A181x_c <= A181x;
			A182x_c <= A182x;
			A183x_c <= A183x;
			A184x_c <= A184x;
			A185x_c <= A185x;
			A186x_c <= A186x;
			sumout<={sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x[15],sum0x}+{sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x[15],sum1x}+{sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x[15],sum2x}+{sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x[15],sum3x}+{sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x[15],sum4x}+{sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x[15],sum5x}+{sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x[15],sum6x}+{sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x[15],sum7x}+{sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x[15],sum8x}+{sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x[15],sum9x}+{sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x[15],sum10x}+{sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x[15],sum11x}+{sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x[15],sum12x}+{sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x[15],sum13x}+{sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x[15],sum14x}+{sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x[15],sum15x}+{sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x[15],sum16x}+{sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x[15],sum17x}+{sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x[15],sum18x}+{sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x[15],sum19x}+{sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x[15],sum20x}+{sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x[15],sum21x}+{sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x[15],sum22x}+{sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x[15],sum23x}+{sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x[15],sum24x}+{sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x[15],sum25x}+{sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x[15],sum26x}+{sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x[15],sum27x}+{sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x[15],sum28x}+{sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x[15],sum29x}+{sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x[15],sum30x}+{sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x[15],sum31x}+{sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x[15],sum32x}+{sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x[15],sum33x}+{sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x[15],sum34x}+{sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x[15],sum35x}+{sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x[15],sum36x}+{sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x[15],sum37x}+{sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x[15],sum38x}+{sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x[15],sum39x}+{sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x[15],sum40x}+{sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x[15],sum41x}+{sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x[15],sum42x}+{sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x[15],sum43x}+{sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x[15],sum44x}+{sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x[15],sum45x}+{sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x[15],sum46x}+{sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x[15],sum47x}+{sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x[15],sum48x}+{sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x[15],sum49x}+{sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x[15],sum50x}+{sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x[15],sum51x}+{sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x[15],sum52x}+{sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x[15],sum53x}+{sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x[15],sum54x}+{sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x[15],sum55x}+{sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x[15],sum56x}+{sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x[15],sum57x}+{sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x[15],sum58x}+{sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x[15],sum59x}+{sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x[15],sum60x}+{sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x[15],sum61x}+{sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x[15],sum62x}+{sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x[15],sum63x}+{sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x[15],sum64x}+{sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x[15],sum65x}+{sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x[15],sum66x}+{sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x[15],sum67x}+{sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x[15],sum68x}+{sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x[15],sum69x}+{sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x[15],sum70x}+{sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x[15],sum71x}+{sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x[15],sum72x}+{sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x[15],sum73x}+{sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x[15],sum74x}+{sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x[15],sum75x}+{sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x[15],sum76x}+{sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x[15],sum77x}+{sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x[15],sum78x}+{sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x[15],sum79x}+{sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x[15],sum80x}+{sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x[15],sum81x}+{sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x[15],sum82x}+{sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x[15],sum83x}+{sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x[15],sum84x}+{sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x[15],sum85x}+{sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x[15],sum86x}+{sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x[15],sum87x}+{sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x[15],sum88x}+{sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x[15],sum89x}+{sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x[15],sum90x}+{sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x[15],sum91x}+{sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x[15],sum92x}+{sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x[15],sum93x}+{sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x[15],sum94x}+{sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x[15],sum95x}+{sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x[15],sum96x}+{sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x[15],sum97x}+{sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x[15],sum98x}+{sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x[15],sum99x}+{sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x[15],sum100x}+{sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x[15],sum101x}+{sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x[15],sum102x}+{sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x[15],sum103x}+{sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x[15],sum104x}+{sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x[15],sum105x}+{sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x[15],sum106x}+{sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x[15],sum107x}+{sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x[15],sum108x}+{sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x[15],sum109x}+{sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x[15],sum110x}+{sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x[15],sum111x}+{sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x[15],sum112x}+{sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x[15],sum113x}+{sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x[15],sum114x}+{sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x[15],sum115x}+{sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x[15],sum116x}+{sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x[15],sum117x}+{sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x[15],sum118x}+{sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x[15],sum119x}+{sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x[15],sum120x}+{sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x[15],sum121x}+{sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x[15],sum122x}+{sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x[15],sum123x}+{sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x[15],sum124x}+{sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x[15],sum125x}+{sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x[15],sum126x}+{sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x[15],sum127x}+{sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x[15],sum128x}+{sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x[15],sum129x}+{sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x[15],sum130x}+{sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x[15],sum131x}+{sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x[15],sum132x}+{sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x[15],sum133x}+{sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x[15],sum134x}+{sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x[15],sum135x}+{sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x[15],sum136x}+{sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x[15],sum137x}+{sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x[15],sum138x}+{sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x[15],sum139x}+{sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x[15],sum140x}+{sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x[15],sum141x}+{sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x[15],sum142x}+{sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x[15],sum143x}+{sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x[15],sum144x}+{sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x[15],sum145x}+{sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x[15],sum146x}+{sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x[15],sum147x}+{sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x[15],sum148x}+{sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x[15],sum149x}+{sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x[15],sum150x}+{sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x[15],sum151x}+{sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x[15],sum152x}+{sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x[15],sum153x}+{sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x[15],sum154x}+{sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x[15],sum155x}+{sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x[15],sum156x}+{sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x[15],sum157x}+{sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x[15],sum158x}+{sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x[15],sum159x}+{sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x[15],sum160x}+{sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x[15],sum161x}+{sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x[15],sum162x}+{sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x[15],sum163x}+{sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x[15],sum164x}+{sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x[15],sum165x}+{sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x[15],sum166x}+{sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x[15],sum167x}+{sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x[15],sum168x}+{sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x[15],sum169x}+{sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x[15],sum170x}+{sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x[15],sum171x}+{sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x[15],sum172x}+{sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x[15],sum173x}+{sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x[15],sum174x}+{sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x[15],sum175x}+{sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x[15],sum176x}+{sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x[15],sum177x}+{sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x[15],sum178x}+{sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x[15],sum179x}+{sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x[15],sum180x}+{sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x[15],sum181x}+{sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x[15],sum182x}+{sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x[15],sum183x}+{sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x[15],sum184x}+{sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x[15],sum185x}+{sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x[15],sum186x}+{B0x[15],B0x[15],B0x[15],B0x[15],B0x[15],B0x[15],B0x[15],B0x};

			if(sumout[22]==0)
				begin
				if(sumout[21:13]!=9'b0)
					N3x<=8'd127;
				else
					begin
					if(sumout[5]==1)
						N3x<=sumout[13:6]+8'd1;
					else
						N3x<=sumout[13:6];
					end
				end
			else
				N3x<=8'd0;
			end
		end
endmodule
