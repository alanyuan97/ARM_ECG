module rom_input(EN, clk, I0x, I1x, I2x, I3x, I4x, I5x, I6x, I7x, I8x, I9x, I10x, I11x, I12x, I13x, I14x, I15x, I16x, I17x, I18x, I19x, I20x, I21x, I22x, I23x, I24x, I25x, I26x, I27x, I28x, I29x, I30x, I31x, I32x, I33x, I34x, I35x, I36x, I37x, I38x, I39x, I40x, I41x, I42x, I43x, I44x, I45x, I46x, I47x, I48x, I49x, I50x, I51x, I52x, I53x, I54x, I55x, I56x, I57x, I58x, I59x, I60x, I61x, I62x, I63x, I64x, I65x, I66x, I67x, I68x, I69x, I70x, I71x, I72x, I73x, I74x);
	input EN, clk;
	output reg [7:0] I0x, I1x, I2x, I3x, I4x, I5x, I6x, I7x, I8x, I9x, I10x, I11x, I12x, I13x, I14x, I15x, I16x, I17x, I18x, I19x, I20x, I21x, I22x, I23x, I24x, I25x, I26x, I27x, I28x, I29x, I30x, I31x, I32x, I33x, I34x, I35x, I36x, I37x, I38x, I39x, I40x, I41x, I42x, I43x, I44x, I45x, I46x, I47x, I48x, I49x, I50x, I51x, I52x, I53x, I54x, I55x, I56x, I57x, I58x, I59x, I60x, I61x, I62x, I63x, I64x, I65x, I66x, I67x, I68x, I69x, I70x, I71x, I72x, I73x, I74x;
always@(posedge clk)
	begin
	I0x = 8'd45;
	I1x = 8'd35;
	I2x = -8'd3;
	I3x = 8'd9;
	I4x = 8'd4;
	I5x = 8'd9;
	I6x = 8'd6;
	I7x = 8'd9;
	I8x = 8'd8;
	I9x = 8'd12;
	I10x = 8'd11;
	I11x = 8'd16;
	I12x = 8'd17;
	I13x = 8'd23;
	I14x = 8'd22;
	I15x = 8'd23;
	I16x = 8'd16;
	I17x = 8'd12;
	I18x = 8'd8;
	I19x = 8'd8;
	I20x = 8'd7;
	I21x = 8'd8;
	I22x = 8'd7;
	I23x = 8'd8;
	I24x = 8'd7;
	I25x = 8'd8;
	I26x = 8'd7;
	I27x = 8'd8;
	I28x = 8'd6;
	I29x = 8'd7;
	I30x = 8'd6;
	I31x = 8'd7;
	I32x = 8'd6;
	I33x = 8'd7;
	I34x = 8'd6;
	I35x = 8'd6;
	I36x = 8'd5;
	I37x = 8'd7;
	I38x = 8'd5;
	I39x = 8'd7;
	I40x = 8'd6;
	I41x = 8'd7;
	I42x = 8'd5;
	I43x = 8'd9;
	I44x = 8'd11;
	I45x = 8'd15;
	I46x = 8'd12;
	I47x = 8'd10;
	I48x = 8'd4;
	I49x = 8'd7;
	I50x = 8'd0;
	I51x = 8'd26;
	I52x = 8'd60;
	I53x = 8'd11;
	I54x = 8'd5;
	I55x = 8'd8;
	I56x = 8'd8;
	I57x = 8'd9;
	I58x = 8'd9;
	I59x = 8'd11;
	I60x = 8'd11;
	I61x = 8'd13;
	I62x = 8'd1;
	I63x = 8'd0;
	I64x = 8'd0;
	I65x = 8'd1;
	I66x = -8'd1;
	I67x = 8'd1;
	I68x = -8'd1;
	I69x = 8'd1;
	I70x = -8'd1;
	I71x = 8'd2;
	I72x = -8'd2;
	I73x = 8'd3;
	I74x = -8'd6;
	end
endmodule
