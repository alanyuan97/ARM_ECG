module layer_4(reset,clk,N1x,N2x,N3x,N4x,N5x,N6x,N7x,N8x,N9x,N10x,N11x,N12x,N13x,N14x,N15x,N16x,N17x,N18x,N19x,N20x,N21x,N22x,N23x,N24x,N25x,N26x,N27x,N28x,N29x,N30x,R0x,R1x,R2x,R3x,R4x,R5x,R6x,R7x,R8x,R9x,R10x,R11x,R12x,R13x,R14x);
	input reset, clk; 
	output [23:0] N1x,N2x,N3x,N4x,N5x,N6x,N7x,N8x,N9x,N10x,N11x,N12x,N13x,N14x,N15x,N16x,N17x,N18x,N19x,N20x,N21x,N22x,N23x,N24x,N25x,N26x,N27x,N28x,N29x,N30x;
	input [23:0] R0x,R1x,R2x,R3x,R4x,R5x,R6x,R7x,R8x,R9x,R10x,R11x,R12x,R13x,R14x;

	node4_1 node4_1( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N1x(N1x) 
	); 
	node4_2 node4_2( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N2x(N2x) 
	); 
	node4_3 node4_3( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N3x(N3x) 
	); 
	node4_4 node4_4( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N4x(N4x) 
	); 
	node4_5 node4_5( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N5x(N5x) 
	); 
	node4_6 node4_6( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N6x(N6x) 
	); 
	node4_7 node4_7( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N7x(N7x) 
	); 
	node4_8 node4_8( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N8x(N8x) 
	); 
	node4_9 node4_9( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N9x(N9x) 
	); 
	node4_10 node4_10( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N10x(N10x) 
	); 
	node4_11 node4_11( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N11x(N11x) 
	); 
	node4_12 node4_12( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N12x(N12x) 
	); 
	node4_13 node4_13( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N13x(N13x) 
	); 
	node4_14 node4_14( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N14x(N14x) 
	); 
	node4_15 node4_15( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N15x(N15x) 
	); 
	node4_16 node4_16( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N16x(N16x) 
	); 
	node4_17 node4_17( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N17x(N17x) 
	); 
	node4_18 node4_18( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N18x(N18x) 
	); 
	node4_19 node4_19( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N19x(N19x) 
	); 
	node4_20 node4_20( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N20x(N20x) 
	); 
	node4_21 node4_21( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N21x(N21x) 
	); 
	node4_22 node4_22( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N22x(N22x) 
	); 
	node4_23 node4_23( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N23x(N23x) 
	); 
	node4_24 node4_24( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N24x(N24x) 
	); 
	node4_25 node4_25( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N25x(N25x) 
	); 
	node4_26 node4_26( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N26x(N26x) 
	); 
	node4_27 node4_27( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N27x(N27x) 
	); 
	node4_28 node4_28( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N28x(N28x) 
	); 
	node4_29 node4_29( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N29x(N29x) 
	); 
	node4_30 node4_30( 
		.A0x(R0x), 
		.A1x(R1x), 
		.A2x(R2x), 
		.A3x(R3x), 
		.A4x(R4x), 
		.A5x(R5x), 
		.A6x(R6x), 
		.A7x(R7x), 
		.A8x(R8x), 
		.A9x(R9x), 
		.A10x(R10x), 
		.A11x(R11x), 
		.A12x(R12x), 
		.A13x(R13x), 
		.A14x(R14x), 
		.clk(clk), 
		.reset(reset), 
		.N30x(N30x) 
	); 
endmodule
