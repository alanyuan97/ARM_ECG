module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [7:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [7:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = -30;
	I1x = 63;
	I2x = 46;
	I3x = -26;
	I4x = -23;
	I5x = 47;
	I6x = -24;
	I7x = 39;
	I8x = 47;
	I9x = 55;
	I10x = 21;
	I11x = 17;
	I12x = -51;
	I13x = -61;
	I14x = -25;
	I15x = 10;
	I16x = 1;
	I17x = -33;
	I18x = -24;
	I19x = -56;
	I20x = -46;
	I21x = 3;
	I22x = 42;
	I23x = -59;
	I24x = -2;
	I25x = -38;
	I26x = -60;
	I27x = -1;
	I28x = 24;
	I29x = -38;
	I30x = -59;
	I31x = 14;
	I32x = 51;
	I33x = 46;
	I34x = 0;
	I35x = 21;
	I36x = -20;
	I37x = 48;
	I38x = 0;
	I39x = 49;
	I40x = -42;
	I41x = -34;
	I42x = -20;
	I43x = 46;
	I44x = -35;
	I45x = 35;
	I46x = 2;
	I47x = -26;
	I48x = 48;
	I49x = -18;
	I50x = -20;
	I51x = -6;
	I52x = 27;
	I53x = -7;
	I54x = -50;
	I55x = -42;
	I56x = -27;
	I57x = -11;
	I58x = -10;
	I59x = -47;
	I60x = -38;
	I61x = 14;
	I62x = 60;
	I63x = 6;
	I64x = -23;
	I65x = -8;
	I66x = 39;
	I67x = -25;
	I68x = 7;
	I69x = 24;
	I70x = -51;
	I71x = 47;
	I72x = 3;
	I73x = -5;
	I74x = 60;
	I75x = -28;
	I76x = 18;
	I77x = -25;
	I78x = -24;
	I79x = 54;
	I80x = -45;
	I81x = 0;
	I82x = 12;
	I83x = 10;
	I84x = 31;
	I85x = 54;
	I86x = 52;
	I87x = 41;
	I88x = 17;
	I89x = -58;
	I90x = 26;
	I91x = -17;
	I92x = -37;
	I93x = 15;
	I94x = -39;
	I95x = 22;
	I96x = -43;
	I97x = -18;
	I98x = -14;
	I99x = -16;
	I100x = -39;
	I101x = -56;
	I102x = 55;
	I103x = -51;
	I104x = 27;
	I105x = 16;
	I106x = 18;
	I107x = 4;
	I108x = 42;
	I109x = -55;
	I110x = -63;
	I111x = -3;
	I112x = 4;
	I113x = -19;
	I114x = -33;
	I115x = 0;
	I116x = -29;
	I117x = -20;
	I118x = -55;
	I119x = 55;
	I120x = 5;
	I121x = 36;
	I122x = 22;
	I123x = 17;
	I124x = -63;
	I125x = 21;
	I126x = 31;
	I127x = 2;
	I128x = -23;
	I129x = -60;
	I130x = -15;
	I131x = -16;
	I132x = -58;
	I133x = -20;
	I134x = 15;
	I135x = -4;
	I136x = 32;
	I137x = -43;
	I138x = -4;
	I139x = -42;
	I140x = -30;
	I141x = 46;
	I142x = 34;
	I143x = -55;
	I144x = -13;
	I145x = 59;
	I146x = 41;
	I147x = 52;
	I148x = -27;
	I149x = -27;
	I150x = -41;
	I151x = 36;
	I152x = -19;
	I153x = 38;
	I154x = 5;
	I155x = -8;
	I156x = 57;
	I157x = 49;
	I158x = -43;
	I159x = -63;
	I160x = 30;
	I161x = -12;
	I162x = 15;
	I163x = 19;
	I164x = -12;
	I165x = 12;
	I166x = -29;
	I167x = 53;
	I168x = -8;
	I169x = -42;
	I170x = -57;
	I171x = 17;
	I172x = 36;
	I173x = -32;
	I174x = -42;
	I175x = 36;
	I176x = -46;
	I177x = -53;
	I178x = -3;
	I179x = 25;
	I180x = 0;
	I181x = 51;
	I182x = 18;
	I183x = -31;
	I184x = -44;
	I185x = 22;
	I186x = -21;
	end
endmodule
[1.16694046 0.         0.32390326 0.         0.96730607] 

 [74, 0, 20, 0, 61] 

 ['01001010', '00000000', '00010100', '00000000', '00111101']
