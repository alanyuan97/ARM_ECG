module rom_ary(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 32'b00111111011011011001011111111011;
	I1x = 32'b00111110111101111110010011111011;
	I2x = 32'b00111110010110101101100110000000;
	I3x = 32'b00000000000000000000000000000000;
	I4x = 32'b00111101001001001101000000001011;
	I5x = 32'b00111101111000000100000011011000;
	I6x = 32'b00111101110000010010111010011011;
	I7x = 32'b00111101111110001001000111100110;
	I8x = 32'b00111101111001000100111001011011;
	I9x = 32'b00111101101101100101111111101010;
	I10x = 32'b00111101110110010111111110101010;
	I11x = 32'b00111101101001100010100111100001;
	I12x = 32'b00111110000000011011000001001100;
	I13x = 32'b00111101111100011101000010111000;
	I14x = 32'b00111101111101001000010001100100;
	I15x = 32'b00111110000001010001000011100011;
	I16x = 32'b00111110001101010000011000010100;
	I17x = 32'b00111110000110001010011110000100;
	I18x = 32'b00111101111110001001000111100110;
	I19x = 32'b00111110010000101000100001110001;
	I20x = 32'b00111110000011110011001010101001;
	I21x = 32'b00111110000001111100010010001111;
	I22x = 32'b00111110001101100101111111101010;
	I23x = 32'b00111110000001100110101010111001;
	I24x = 32'b00111110010000001000000110110000;
	I25x = 32'b00111110001001000010001100100000;
	I26x = 32'b00111110010001010011110000011110;
	I27x = 32'b00111110011101001000010001100100;
	I28x = 32'b00111110011010011011010110110011;
	I29x = 32'b00111110011110111111001001111110;
	I30x = 32'b00111110100000001010110011101011;
	I31x = 32'b00111110101001011101001101101011;
	I32x = 32'b00111110110000101101111011100111;
	I33x = 32'b00111110101101111011100111000001;
	I34x = 32'b00111110111010111011110001110100;
	I35x = 32'b00111110110110101000001100001010;
	I36x = 32'b00111110111101111000111010000110;
	I37x = 32'b00111110110111111001001111101101;
	I38x = 32'b00111110110010000100011000111111;
	I39x = 32'b00111110101101100000100101110101;
	I40x = 32'b00111110100100101110100110110110;
	I41x = 32'b00111110100011010010101111101000;
	I42x = 32'b00111110100110101010111001000101;
	I43x = 32'b00111110011011010001011001001010;
	I44x = 32'b00111110011011100111000000100000;
	I45x = 32'b00111110011000011001101010101110;
	I46x = 32'b00111110011000000100000011011000;
	I47x = 32'b00111110010100101011111001111011;
	I48x = 32'b00111110000101010100011011101100;
	I49x = 32'b00111110001111111101010011000101;
	I50x = 32'b00111110010110000010010111010011;
	I51x = 32'b00111110010001110100001011011111;
	I52x = 32'b00111110010111101110011100000010;
	I53x = 32'b00111110001011001110101100010000;
	I54x = 32'b00111110011001001111101101000110;
	I55x = 32'b00111110011001100101010100011100;
	I56x = 32'b00111110010000011101101110000110;
	I57x = 32'b00111110011010010000100011001000;
	I58x = 32'b00111110010011010101011100100010;
	I59x = 32'b00111110011000101111010010000100;
	I60x = 32'b00111110011101011101111000111010;
	I61x = 32'b00111110010101000001100001010001;
	I62x = 32'b00111110010101100001111100010010;
	I63x = 32'b00111110001100000100101110100111;
	I64x = 32'b00111110011001011010100000110001;
	I65x = 32'b00111110011000001110110111000011;
	I66x = 32'b00111110011010100110001010011110;
	I67x = 32'b00111110100000101011001110101100;
	I68x = 32'b00111110001011111001111010111100;
	I69x = 32'b00111110010001111110111111001010;
	I70x = 32'b00111110010110101101100110000000;
	I71x = 32'b00111110010101110111100011101000;
	I72x = 32'b00111110010011001010101000110111;
	I73x = 32'b00111110001111110010011111011010;
	I74x = 32'b00111110010100101011111001111011;
	I75x = 32'b00111110010111111001001111101101;
	I76x = 32'b00111110010100001011011110111010;
	I77x = 32'b00111110011011011100001100110101;
	I78x = 32'b00111110000011101000010110111110;
	I79x = 32'b00111110010101001100010100111100;
	I80x = 32'b00111110100000010000001101100001;
	I81x = 32'b00111110010011001010101000110111;
	I82x = 32'b00111110010110001101001010111110;
	I83x = 32'b00111110000110010101010001101111;
	I84x = 32'b00111110001011000011111000100100;
	I85x = 32'b00111110001100011010010101111101;
	I86x = 32'b00111110001011101111000111010001;
	I87x = 32'b00111110010100010110010010100101;
	I88x = 32'b00111101111101011101111000111010;
	I89x = 32'b00111110001111010010000100011001;
	I90x = 32'b00111110000110101010111001000101;
	I91x = 32'b00111110001111000111010000101110;
	I92x = 32'b00111110001111000111010000101110;
	I93x = 32'b00111110000110100000000101011010;
	I94x = 32'b00111110001100100101001001101000;
	I95x = 32'b00111110011000000100000011011000;
	I96x = 32'b00111110001010111001000100111001;
	I97x = 32'b00111110010010010100100110100000;
	I98x = 32'b00111110010111001110000001000001;
	I99x = 32'b00111110100000000000000000000000;
	I100x = 32'b00111110100001110001011110100100;
	I101x = 32'b00111110100111001011010100000110;
	I102x = 32'b00111110100101001001101000000001;
	I103x = 32'b00111110100011101000010110111110;
	I104x = 32'b00111110100111010110000111110001;
	I105x = 32'b00111110100110100000000101011010;
	I106x = 32'b00111110100011100010111101001000;
	I107x = 32'b00111110100101110100110110101110;
	I108x = 32'b00111110011011000110100101011111;
	I109x = 32'b00111110011010010000100011001000;
	I110x = 32'b00111110001110000110011010101100;
	I111x = 32'b00111110001110000110011010101100;
	I112x = 32'b00111110010000111110001001001000;
	I113x = 32'b00111110000111100000111011011100;
	I114x = 32'b00111110011100111101011101111001;
	I115x = 32'b00111110010100110110101101100110;
	I116x = 32'b00111110001101111011100111000001;
	I117x = 32'b00111110001010101110010001001110;
	I118x = 32'b00111110101001111000001110110111;
	I119x = 32'b00111111000111010011011010110110;
	I120x = 32'b00111111100000000000000000000000;
	I121x = 32'b00111111000001101001010111110100;
	I122x = 32'b00111110100000010000001101100001;
	I123x = 32'b00111101010110101101100110000000;
	I124x = 32'b00111110000111100000111011011100;
	I125x = 32'b00111110001111100111101011101111;
	I126x = 32'b00111110001111100111101011101111;
	I127x = 32'b00111110010100010110010010100101;
	I128x = 32'b00111110001110110001101001011000;
	I129x = 32'b00111110001011101111000111010001;
	I130x = 32'b00111110001011101111000111010001;
	I131x = 32'b00111110000111110110100010110010;
	I132x = 32'b00111110001011101111000111010001;
	I133x = 32'b00111110001111011100111000000100;
	I134x = 32'b00111110011101011101111000111010;
	I135x = 32'b00111110001110111100011101000011;
	I136x = 32'b00111110001100001111100010010010;
	I137x = 32'b00111110000111100000111011011100;
	I138x = 32'b00111110000111110110100010110010;
	I139x = 32'b00111110010111001110000001000001;
	I140x = 32'b00111110010001110100001011011111;
	I141x = 32'b00000000000000000000000000000000;
	I142x = 32'b00000000000000000000000000000000;
	I143x = 32'b00000000000000000000000000000000;
	I144x = 32'b00000000000000000000000000000000;
	I145x = 32'b00000000000000000000000000000000;
	I146x = 32'b00000000000000000000000000000000;
	I147x = 32'b00000000000000000000000000000000;
	I148x = 32'b00000000000000000000000000000000;
	I149x = 32'b00000000000000000000000000000000;
	I150x = 32'b00000000000000000000000000000000;
	I151x = 32'b00000000000000000000000000000000;
	I152x = 32'b00000000000000000000000000000000;
	I153x = 32'b00000000000000000000000000000000;
	I154x = 32'b00000000000000000000000000000000;
	I155x = 32'b00000000000000000000000000000000;
	I156x = 32'b00000000000000000000000000000000;
	I157x = 32'b00000000000000000000000000000000;
	I158x = 32'b00000000000000000000000000000000;
	I159x = 32'b00000000000000000000000000000000;
	I160x = 32'b00000000000000000000000000000000;
	I161x = 32'b00000000000000000000000000000000;
	I162x = 32'b00000000000000000000000000000000;
	I163x = 32'b00000000000000000000000000000000;
	I164x = 32'b00000000000000000000000000000000;
	I165x = 32'b00000000000000000000000000000000;
	I166x = 32'b00000000000000000000000000000000;
	I167x = 32'b00000000000000000000000000000000;
	I168x = 32'b00000000000000000000000000000000;
	I169x = 32'b00000000000000000000000000000000;
	I170x = 32'b00000000000000000000000000000000;
	I171x = 32'b00000000000000000000000000000000;
	I172x = 32'b00000000000000000000000000000000;
	I173x = 32'b00000000000000000000000000000000;
	I174x = 32'b00000000000000000000000000000000;
	I175x = 32'b00000000000000000000000000000000;
	I176x = 32'b00000000000000000000000000000000;
	I177x = 32'b00000000000000000000000000000000;
	I178x = 32'b00000000000000000000000000000000;
	I179x = 32'b00000000000000000000000000000000;
	I180x = 32'b00000000000000000000000000000000;
	I181x = 32'b00000000000000000000000000000000;
	I182x = 32'b00000000000000000000000000000000;
	I183x = 32'b00000000000000000000000000000000;
	I184x = 32'b00000000000000000000000000000000;
	I185x = 32'b00000000000000000000000000000000;
	I186x = 32'b00000000000000000000000000000000;
	end
endmodule