module rom_rand1(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 274;   
	I1x = -819;
	I2x = -229;
	I3x = 194;
	I4x = 392;
	I5x = -26;
	I6x = -49;
	I7x = 364;
	I8x = 42;
	I9x = -475;
	I10x = -593;
	I11x = 479;
	I12x = 463;
	I13x = -946;
	I14x = -1016;
	I15x = 255;
	I16x = 889;
	I17x = -783;
	I18x = 789;
	I19x = -698;
	I20x = -27;
	I21x = -614;
	I22x = 1018;
	I23x = 651;
	I24x = -730;
	I25x = 831;
	I26x = 179;
	I27x = -314;
	I28x = 195;
	I29x = -497;
	I30x = 639;
	I31x = 832;
	I32x = 338;
	I33x = -22;
	I34x = 158;
	I35x = 149;
	I36x = -450;
	I37x = 89;
	I38x = -381;
	I39x = 659;
	I40x = 122;
	I41x = 141;
	I42x = 365;
	I43x = 519;
	I44x = 860;
	I45x = -17;
	I46x = 694;
	I47x = 888;
	I48x = -596;
	I49x = 735;
	I50x = -287;
	I51x = -141;
	I52x = 243;
	I53x = 897;
	I54x = 925;
	I55x = -641;
	I56x = -672;
	I57x = -491;
	I58x = -230;
	I59x = -896;
	I60x = 82;
	I61x = -610;
	I62x = -216;
	I63x = 33;
	I64x = 725;
	I65x = -527;
	I66x = -1009;
	I67x = 483;
	I68x = 276;
	I69x = -922;
	I70x = -92;
	I71x = -35;
	I72x = -34;
	I73x = 788;
	I74x = -541;
	I75x = 60;
	I76x = 893;
	I77x = -705;
	I78x = 173;
	I79x = -512;
	I80x = -336;
	I81x = 719;
	I82x = 850;
	I83x = 538;
	I84x = -556;
	I85x = -312;
	I86x = -873;
	I87x = -459;
	I88x = 374;
	I89x = 646;
	I90x = -42;
	I91x = -236;
	I92x = -551;
	I93x = 114;
	I94x = -635;
	I95x = -231;
	I96x = -97;
	I97x = 607;
	I98x = -758;
	I99x = 814;
	I100x = 751;
	I101x = 92;
	I102x = 25;
	I103x = 847;
	I104x = 86;
	I105x = -355;
	I106x = 667;
	I107x = 6;
	I108x = 574;
	I109x = -134;
	I110x = 952;
	I111x = 623;
	I112x = -692;
	I113x = 860;
	I114x = -630;
	I115x = 273;
	I116x = 845;
	I117x = -917;
	I118x = 95;
	I119x = 485;
	I120x = 469;
	I121x = 645;
	I122x = 628;
	I123x = 331;
	I124x = -617;
	I125x = -928;
	I126x = -230;
	I127x = -756;
	I128x = 500;
	I129x = 910;
	I130x = -606;
	I131x = -355;
	I132x = -629;
	I133x = -990;
	I134x = 29;
	I135x = -207;
	I136x = 700;
	I137x = 352;
	I138x = 223;
	I139x = 277;
	I140x = 500;
	I141x = 767;
	I142x = -327;
	I143x = -361;
	I144x = 872;
	I145x = 156;
	I146x = 324;
	I147x = -741;
	I148x = 338;
	I149x = -44;
	I150x = -608;
	I151x = -953;
	I152x = -107;
	I153x = -222;
	I154x = -738;
	I155x = 774;
	I156x = 740;
	I157x = -83;
	I158x = 752;
	I159x = 333;
	I160x = 308;
	I161x = -182;
	I162x = 574;
	I163x = 302;
	I164x = 561;
	I165x = 609;
	I166x = 28;
	I167x = 801;
	I168x = -144;
	I169x = 443;
	I170x = -285;
	I171x = 626;
	I172x = -1001;
	I173x = -535;
	I174x = 283;
	I175x = 98;
	I176x = 128;
	I177x = -525;
	I178x = 579;
	I179x = -541;
	I180x = 204;
	I181x = -271;
	I182x = -700;
	I183x = 439;
	I184x = -137;
	I185x = 810;
	I186x = 276;
	end
endmodule