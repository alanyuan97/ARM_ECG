module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 1024;
	I1x = 822;
	I2x = 228;
	I3x = 20;
	I4x = 101;
	I5x = 136;
	I6x = 106;
	I7x = 130;
	I8x = 145;
	I9x = 128;
	I10x = 176;
	I11x = 159;
	I12x = 173;
	I13x = 171;
	I14x = 152;
	I15x = 190;
	I16x = 175;
	I17x = 189;
	I18x = 187;
	I19x = 171;
	I20x = 208;
	I21x = 191;
	I22x = 201;
	I23x = 206;
	I24x = 187;
	I25x = 233;
	I26x = 229;
	I27x = 241;
	I28x = 246;
	I29x = 227;
	I30x = 275;
	I31x = 260;
	I32x = 261;
	I33x = 257;
	I34x = 234;
	I35x = 268;
	I36x = 241;
	I37x = 237;
	I38x = 224;
	I39x = 192;
	I40x = 227;
	I41x = 215;
	I42x = 214;
	I43x = 212;
	I44x = 180;
	I45x = 222;
	I46x = 208;
	I47x = 206;
	I48x = 198;
	I49x = 173;
	I50x = 210;
	I51x = 194;
	I52x = 191;
	I53x = 197;
	I54x = 170;
	I55x = 211;
	I56x = 193;
	I57x = 203;
	I58x = 205;
	I59x = 179;
	I60x = 212;
	I61x = 201;
	I62x = 197;
	I63x = 200;
	I64x = 172;
	I65x = 207;
	I66x = 193;
	I67x = 193;
	I68x = 205;
	I69x = 183;
	I70x = 228;
	I71x = 219;
	I72x = 233;
	I73x = 243;
	I74x = 221;
	I75x = 246;
	I76x = 242;
	I77x = 229;
	I78x = 208;
	I79x = 128;
	I80x = 184;
	I81x = 175;
	I82x = 191;
	I83x = 193;
	I84x = 148;
	I85x = 177;
	I86x = 196;
	I87x = 315;
	I88x = 496;
	I89x = 569;
	I90x = 834;
	I91x = 1016;
	I92x = 614;
	I93x = 129;
	I94x = 0;
	I95x = 127;
	I96x = 94;
	I97x = 102;
	I98x = 121;
	I99x = 107;
	I100x = 141;
	I101x = 135;
	I102x = 147;
	I103x = 157;
	I104x = 128;
	I105x = 155;
	I106x = 151;
	I107x = 155;
	I108x = 176;
	I109x = 0;
	I110x = 0;
	I111x = 0;
	I112x = 0;
	I113x = 0;
	I114x = 0;
	I115x = 0;
	I116x = 0;
	I117x = 0;
	I118x = 0;
	I119x = 0;
	I120x = 0;
	I121x = 0;
	I122x = 0;
	I123x = 0;
	I124x = 0;
	I125x = 0;
	I126x = 0;
	I127x = 0;
	I128x = 0;
	I129x = 0;
	I130x = 0;
	I131x = 0;
	I132x = 0;
	I133x = 0;
	I134x = 0;
	I135x = 0;
	I136x = 0;
	I137x = 0;
	I138x = 0;
	I139x = 0;
	I140x = 0;
	I141x = 0;
	I142x = 0;
	I143x = 0;
	I144x = 0;
	I145x = 0;
	I146x = 0;
	I147x = 0;
	I148x = 0;
	I149x = 0;
	I150x = 0;
	I151x = 0;
	I152x = 0;
	I153x = 0;
	I154x = 0;
	I155x = 0;
	I156x = 0;
	I157x = 0;
	I158x = 0;
	I159x = 0;
	I160x = 0;
	I161x = 0;
	I162x = 0;
	I163x = 0;
	I164x = 0;
	I165x = 0;
	I166x = 0;
	I167x = 0;
	I168x = 0;
	I169x = 0;
	I170x = 0;
	I171x = 0;
	I172x = 0;
	I173x = 0;
	I174x = 0;
	I175x = 0;
	I176x = 0;
	I177x = 0;
	I178x = 0;
	I179x = 0;
	I180x = 0;
	I181x = 0;
	I182x = 0;
	I183x = 0;
	I184x = 0;
	I185x = 0;
	I186x = 0;
	end
endmodule
