module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [31:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 8036;
	I1x = 6291;
	I2x = 3153;
	I3x = 1433;
	I4x = 0;
	I5x = 109;
	I6x = 599;
	I7x = 892;
	I8x = 950;
	I9x = 1081;
	I10x = 1138;
	I11x = 1171;
	I12x = 1236;
	I13x = 1236;
	I14x = 1196;
	I15x = 1294;
	I16x = 1343;
	I17x = 1409;
	I18x = 1449;
	I19x = 1515;
	I20x = 1564;
	I21x = 1654;
	I22x = 1753;
	I23x = 1818;
	I24x = 2048;
	I25x = 2244;
	I26x = 2424;
	I27x = 2596;
	I28x = 2875;
	I29x = 2932;
	I30x = 3121;
	I31x = 3293;
	I32x = 3416;
	I33x = 3424;
	I34x = 3342;
	I35x = 3309;
	I36x = 3063;
	I37x = 2777;
	I38x = 2473;
	I39x = 2203;
	I40x = 1949;
	I41x = 1884;
	I42x = 1720;
	I43x = 1589;
	I44x = 1589;
	I45x = 1507;
	I46x = 1449;
	I47x = 1409;
	I48x = 1433;
	I49x = 1409;
	I50x = 1417;
	I51x = 1417;
	I52x = 1540;
	I53x = 1589;
	I54x = 1507;
	I55x = 1499;
	I56x = 1458;
	I57x = 1507;
	I58x = 1564;
	I59x = 1556;
	I60x = 1523;
	I61x = 1449;
	I62x = 1490;
	I63x = 1400;
	I64x = 1482;
	I65x = 1507;
	I66x = 1449;
	I67x = 1384;
	I68x = 1449;
	I69x = 1523;
	I70x = 1482;
	I71x = 1482;
	I72x = 1515;
	I73x = 1523;
	I74x = 1572;
	I75x = 1540;
	I76x = 1540;
	I77x = 1572;
	I78x = 1531;
	I79x = 1540;
	I80x = 1474;
	I81x = 1613;
	I82x = 1720;
	I83x = 1859;
	I84x = 2031;
	I85x = 2277;
	I86x = 2441;
	I87x = 2629;
	I88x = 2572;
	I89x = 2572;
	I90x = 2220;
	I91x = 2105;
	I92x = 1941;
	I93x = 1572;
	I94x = 1310;
	I95x = 1269;
	I96x = 1294;
	I97x = 1236;
	I98x = 1302;
	I99x = 1236;
	I100x = 1187;
	I101x = 950;
	I102x = 1310;
	I103x = 3399;
	I104x = 6938;
	I105x = 8192;
	I106x = 6283;
	I107x = 3358;
	I108x = 1777;
	I109x = 340;
	I110x = 439;
	I111x = 966;
	I112x = 1245;
	I113x = 1286;
	I114x = 1310;
	I115x = 1335;
	I116x = 1409;
	I117x = 1425;
	I118x = 1474;
	I119x = 1482;
	I120x = 1458;
	I121x = 1433;
	I122x = 1564;
	I123x = 1564;
	I124x = 1671;
	I125x = 1671;
	I126x = 1761;
	I127x = 1892;
	I128x = 1957;
	I129x = 2056;
	I130x = 2179;
	I131x = 2375;
	I132x = 2547;
	I133x = 2711;
	I134x = 2949;
	I135x = 3080;
	I136x = 3194;
	I137x = 3276;
	I138x = 3317;
	I139x = 3334;
	I140x = 3211;
	I141x = 3031;
	I142x = 2785;
	I143x = 2547;
	I144x = 0;
	I145x = 0;
	I146x = 0;
	I147x = 0;
	I148x = 0;
	I149x = 0;
	I150x = 0;
	I151x = 0;
	I152x = 0;
	I153x = 0;
	I154x = 0;
	I155x = 0;
	I156x = 0;
	I157x = 0;
	I158x = 0;
	I159x = 0;
	I160x = 0;
	I161x = 0;
	I162x = 0;
	I163x = 0;
	I164x = 0;
	I165x = 0;
	I166x = 0;
	I167x = 0;
	I168x = 0;
	I169x = 0;
	I170x = 0;
	I171x = 0;
	I172x = 0;
	I173x = 0;
	I174x = 0;
	I175x = 0;
	I176x = 0;
	I177x = 0;
	I178x = 0;
	I179x = 0;
	I180x = 0;
	I181x = 0;
	I182x = 0;
	I183x = 0;
	I184x = 0;
	I185x = 0;
	I186x = 0;
	end
endmodule
