module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [7:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [7:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 16'sb0000000001010111;
	I1x = 16'sb0000000101101100;
	I2x = 16'sb1111111110110100;
	I3x = 16'sb0000000100011001;
	I4x = 16'sb0000001110100011;
	I5x = 16'sb1111110000110010;
	I6x = 16'sb1111110111010010;
	I7x = 16'sb1111111010110111;
	I8x = 16'sb1111110101110111;
	I9x = 16'sb0000001100011101;
	I10x = 16'sb0000001101000011;
	I11x = 16'sb0000000100010111;
	I12x = 16'sb1111111000001001;
	I13x = 16'sb1111111100110001;
	I14x = 16'sb0000001100110001;
	I15x = 16'sb0000000101010000;
	I16x = 16'sb1111111010010000;
	I17x = 16'sb1111111011111110;
	I18x = 16'sb0000001101001111;
	I19x = 16'sb0000001001001000;
	I20x = 16'sb1111110001110000;
	I21x = 16'sb1111110011000100;
	I22x = 16'sb1111110101000010;
	I23x = 16'sb1111111110001101;
	I24x = 16'sb1111110110001101;
	I25x = 16'sb1111111100100100;
	I26x = 16'sb1111111000001111;
	I27x = 16'sb0000001010001011;
	I28x = 16'sb1111111001000111;
	I29x = 16'sb1111111000100001;
	I30x = 16'sb0000001000000101;
	I31x = 16'sb0000000101010010;
	I32x = 16'sb1111110011110000;
	I33x = 16'sb1111110110110101;
	I34x = 16'sb0000000100010111;
	I35x = 16'sb1111111100111111;
	I36x = 16'sb1111111101011000;
	I37x = 16'sb0000001000010101;
	I38x = 16'sb0000001001100111;
	I39x = 16'sb0000001010011111;
	I40x = 16'sb1111110111011100;
	I41x = 16'sb1111110101010001;
	I42x = 16'sb0000000010000101;
	I43x = 16'sb1111111110101010;
	I44x = 16'sb0000000011000111;
	I45x = 16'sb0000000100100010;
	I46x = 16'sb0000000110101101;
	I47x = 16'sb0000000010110100;
	I48x = 16'sb1111110110000101;
	I49x = 16'sb1111110011111010;
	I50x = 16'sb1111110100111111;
	I51x = 16'sb1111110111111010;
	I52x = 16'sb1111110100000010;
	I53x = 16'sb1111111101111111;
	I54x = 16'sb1111110000000111;
	I55x = 16'sb0000000010101011;
	I56x = 16'sb1111110010100110;
	I57x = 16'sb0000000011011101;
	I58x = 16'sb0000000010011100;
	I59x = 16'sb1111111010000101;
	I60x = 16'sb1111110101011100;
	I61x = 16'sb1111111011000001;
	I62x = 16'sb0000001011000110;
	I63x = 16'sb1111110100001110;
	I64x = 16'sb1111111001011011;
	I65x = 16'sb1111111001000010;
	I66x = 16'sb1111111000000010;
	I67x = 16'sb1111111011010101;
	I68x = 16'sb1111111101101110;
	I69x = 16'sb1111111101110001;
	I70x = 16'sb1111110100000101;
	I71x = 16'sb1111110011000000;
	I72x = 16'sb1111111110100010;
	I73x = 16'sb0000001111010110;
	I74x = 16'sb0000001101100000;
	I75x = 16'sb1111111101101100;
	I76x = 16'sb0000001111001100;
	I77x = 16'sb0000000110110010;
	I78x = 16'sb0000001111111111;
	I79x = 16'sb1111111011111110;
	I80x = 16'sb1111111000010011;
	I81x = 16'sb0000000100000111;
	I82x = 16'sb1111110001101111;
	I83x = 16'sb1111110010010000;
	I84x = 16'sb1111110000010111;
	I85x = 16'sb0000000111111011;
	I86x = 16'sb1111110100010010;
	I87x = 16'sb1111110011101101;
	I88x = 16'sb1111111100100101;
	I89x = 16'sb0000001001111010;
	I90x = 16'sb0000000001111011;
	I91x = 16'sb0000000010001011;
	I92x = 16'sb0000001011100110;
	I93x = 16'sb1111111000011111;
	I94x = 16'sb1111110110101111;
	I95x = 16'sb1111110101100100;
	I96x = 16'sb1111111101100011;
	I97x = 16'sb0000001001111010;
	I98x = 16'sb1111111111101100;
	I99x = 16'sb1111110111011111;
	I100x = 16'sb1111110111010110;
	I101x = 16'sb0000000100000111;
	I102x = 16'sb0000000011010110;
	I103x = 16'sb0000001011111000;
	I104x = 16'sb1111111100100010;
	I105x = 16'sb1111111100010011;
	I106x = 16'sb1111110011111011;
	I107x = 16'sb1111110101110100;
	I108x = 16'sb1111110101100010;
	I109x = 16'sb0000001110101010;
	I110x = 16'sb1111111010111111;
	I111x = 16'sb1111110011101110;
	I112x = 16'sb0000001000111011;
	I113x = 16'sb1111111110111011;
	I114x = 16'sb1111110110010010;
	I115x = 16'sb0000001101101010;
	I116x = 16'sb0000000100010100;
	I117x = 16'sb1111111110000110;
	I118x = 16'sb0000001101101111;
	I119x = 16'sb0000000111001100;
	I120x = 16'sb1111111011111101;
	I121x = 16'sb0000001010010111;
	I122x = 16'sb0000000001100111;
	I123x = 16'sb1111111001011110;
	I124x = 16'sb0000000010101011;
	I125x = 16'sb1111110110110011;
	I126x = 16'sb1111111000000000;
	I127x = 16'sb0000000110111001;
	I128x = 16'sb1111111110001110;
	I129x = 16'sb1111111111001111;
	I130x = 16'sb1111110011001011;
	I131x = 16'sb1111111101111010;
	I132x = 16'sb0000001110100011;
	I133x = 16'sb1111110111000110;
	I134x = 16'sb1111110111011010;
	I135x = 16'sb1111111111011100;
	I136x = 16'sb1111110000010011;
	I137x = 16'sb1111111011011011;
	I138x = 16'sb1111110101010010;
	I139x = 16'sb0000000000010000;
	I140x = 16'sb1111111101111100;
	I141x = 16'sb0000001101110101;
	I142x = 16'sb0000000011110001;
	I143x = 16'sb1111110000001111;
	I144x = 16'sb1111111110101011;
	I145x = 16'sb1111111101100000;
	I146x = 16'sb0000000000011101;
	I147x = 16'sb1111110011010010;
	I148x = 16'sb0000001001100000;
	I149x = 16'sb0000000010010110;
	I150x = 16'sb0000000110010100;
	I151x = 16'sb1111110111111000;
	I152x = 16'sb1111111010110011;
	I153x = 16'sb0000001011000000;
	I154x = 16'sb1111111111011001;
	I155x = 16'sb1111110001000100;
	I156x = 16'sb1111111001010111;
	I157x = 16'sb0000000110011011;
	I158x = 16'sb0000001110011110;
	I159x = 16'sb1111111101111110;
	I160x = 16'sb0000001101001101;
	I161x = 16'sb1111111110111111;
	I162x = 16'sb0000001001110010;
	I163x = 16'sb0000000001010000;
	I164x = 16'sb1111111100110110;
	I165x = 16'sb1111111101010100;
	I166x = 16'sb1111110111111101;
	I167x = 16'sb1111111010001011;
	I168x = 16'sb1111110101100001;
	I169x = 16'sb1111110100011011;
	I170x = 16'sb0000000101100111;
	I171x = 16'sb1111111010010110;
	I172x = 16'sb1111111110001000;
	I173x = 16'sb0000000001101001;
	I174x = 16'sb0000000100111001;
	I175x = 16'sb0000001011111110;
	I176x = 16'sb0000000100011001;
	I177x = 16'sb1111110110010001;
	I178x = 16'sb1111110010000000;
	I179x = 16'sb1111110010110101;
	I180x = 16'sb0000000100110111;
	I181x = 16'sb0000001000000010;
	I182x = 16'sb1111110010111000;
	I183x = 16'sb0000000010110110;
	I184x = 16'sb0000001001011100;
	I185x = 16'sb0000000100110001;
	I186x = 16'sb1111111000100110;
	end
endmodule
[0.46984231 0.         1.23969952 2.0304947  0.        ] ["16'sb0000000111100001", "16'sb0000000000000000", "16'sb0000010011110101", "16'sb0000100000011111", "16'sb0000000000000000"]
