module sigmoid_approx()