module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 31;
	I1x = 24;
	I2x = 12;
	I3x = 5;
	I4x = 0;
	I5x = 0;
	I6x = 2;
	I7x = 3;
	I8x = 3;
	I9x = 4;
	I10x = 4;
	I11x = 4;
	I12x = 4;
	I13x = 4;
	I14x = 4;
	I15x = 5;
	I16x = 5;
	I17x = 5;
	I18x = 5;
	I19x = 5;
	I20x = 6;
	I21x = 6;
	I22x = 6;
	I23x = 7;
	I24x = 8;
	I25x = 8;
	I26x = 9;
	I27x = 10;
	I28x = 11;
	I29x = 11;
	I30x = 12;
	I31x = 12;
	I32x = 13;
	I33x = 13;
	I34x = 13;
	I35x = 12;
	I36x = 11;
	I37x = 10;
	I38x = 9;
	I39x = 8;
	I40x = 7;
	I41x = 7;
	I42x = 6;
	I43x = 6;
	I44x = 6;
	I45x = 5;
	I46x = 5;
	I47x = 5;
	I48x = 5;
	I49x = 5;
	I50x = 5;
	I51x = 5;
	I52x = 6;
	I53x = 6;
	I54x = 5;
	I55x = 5;
	I56x = 5;
	I57x = 5;
	I58x = 6;
	I59x = 6;
	I60x = 5;
	I61x = 5;
	I62x = 5;
	I63x = 5;
	I64x = 5;
	I65x = 5;
	I66x = 5;
	I67x = 5;
	I68x = 5;
	I69x = 5;
	I70x = 5;
	I71x = 5;
	I72x = 5;
	I73x = 5;
	I74x = 6;
	I75x = 6;
	I76x = 6;
	I77x = 6;
	I78x = 5;
	I79x = 6;
	I80x = 5;
	I81x = 6;
	I82x = 6;
	I83x = 7;
	I84x = 7;
	I85x = 8;
	I86x = 9;
	I87x = 10;
	I88x = 10;
	I89x = 10;
	I90x = 8;
	I91x = 8;
	I92x = 7;
	I93x = 6;
	I94x = 5;
	I95x = 4;
	I96x = 5;
	I97x = 4;
	I98x = 5;
	I99x = 4;
	I100x = 4;
	I101x = 3;
	I102x = 5;
	I103x = 13;
	I104x = 27;
	I105x = 32;
	I106x = 24;
	I107x = 13;
	I108x = 6;
	I109x = 1;
	I110x = 1;
	I111x = 3;
	I112x = 4;
	I113x = 5;
	I114x = 5;
	I115x = 5;
	I116x = 5;
	I117x = 5;
	I118x = 5;
	I119x = 5;
	I120x = 5;
	I121x = 5;
	I122x = 6;
	I123x = 6;
	I124x = 6;
	I125x = 6;
	I126x = 6;
	I127x = 7;
	I128x = 7;
	I129x = 8;
	I130x = 8;
	I131x = 9;
	I132x = 9;
	I133x = 10;
	I134x = 11;
	I135x = 12;
	I136x = 12;
	I137x = 12;
	I138x = 12;
	I139x = 13;
	I140x = 12;
	I141x = 11;
	I142x = 10;
	I143x = 9;
	I144x = 0;
	I145x = 0;
	I146x = 0;
	I147x = 0;
	I148x = 0;
	I149x = 0;
	I150x = 0;
	I151x = 0;
	I152x = 0;
	I153x = 0;
	I154x = 0;
	I155x = 0;
	I156x = 0;
	I157x = 0;
	I158x = 0;
	I159x = 0;
	I160x = 0;
	I161x = 0;
	I162x = 0;
	I163x = 0;
	I164x = 0;
	I165x = 0;
	I166x = 0;
	I167x = 0;
	I168x = 0;
	I169x = 0;
	I170x = 0;
	I171x = 0;
	I172x = 0;
	I173x = 0;
	I174x = 0;
	I175x = 0;
	I176x = 0;
	I177x = 0;
	I178x = 0;
	I179x = 0;
	I180x = 0;
	I181x = 0;
	I182x = 0;
	I183x = 0;
	I184x = 0;
	I185x = 0;
	I186x = 0;
	end
endmodule
