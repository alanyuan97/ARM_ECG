module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = -4425;
	I1x = -2387;
	I2x = 3029;
	I3x = -7163;
	I4x = 7977;
	I5x = 353;
	I6x = 5078;
	I7x = -2826;
	I8x = 4335;
	I9x = -126;
	I10x = -3120;
	I11x = -1204;
	I12x = 386;
	I13x = 4529;
	I14x = 1969;
	I15x = 4683;
	I16x = 468;
	I17x = 2894;
	I18x = 1656;
	I19x = -2835;
	I20x = -4994;
	I21x = 1057;
	I22x = -961;
	I23x = -4640;
	I24x = -5445;
	I25x = 7218;
	I26x = -1018;
	I27x = -8086;
	I28x = -5920;
	I29x = 5205;
	I30x = 821;
	I31x = 4225;
	I32x = -4737;
	I33x = 8123;
	I34x = -3121;
	I35x = -1746;
	I36x = -3455;
	I37x = -4555;
	I38x = -3982;
	I39x = -6582;
	I40x = 5755;
	I41x = -5414;
	I42x = 5446;
	I43x = 3967;
	I44x = -7247;
	I45x = -7393;
	I46x = 775;
	I47x = -6020;
	I48x = -7452;
	I49x = 5663;
	I50x = -5212;
	I51x = -962;
	I52x = -1536;
	I53x = 572;
	I54x = 7108;
	I55x = -7414;
	I56x = 5384;
	I57x = 7061;
	I58x = 2084;
	I59x = 5256;
	I60x = -6854;
	I61x = 6781;
	I62x = 7043;
	I63x = -3810;
	I64x = 7338;
	I65x = -6520;
	I66x = 7214;
	I67x = -494;
	I68x = 1196;
	I69x = -4942;
	I70x = 4744;
	I71x = -1825;
	I72x = -2710;
	I73x = 7042;
	I74x = 1256;
	I75x = 5430;
	I76x = -7352;
	I77x = -1780;
	I78x = 1579;
	I79x = 6287;
	I80x = 1421;
	I81x = 4198;
	I82x = -3116;
	I83x = -3397;
	I84x = 507;
	I85x = -4356;
	I86x = -121;
	I87x = 2438;
	I88x = -3327;
	I89x = -2350;
	I90x = -5642;
	I91x = -7229;
	I92x = 3321;
	I93x = 7546;
	I94x = -5695;
	I95x = -2028;
	I96x = -297;
	I97x = 2181;
	I98x = -4880;
	I99x = 1734;
	I100x = -7048;
	I101x = 4739;
	I102x = -7355;
	I103x = 1859;
	I104x = -479;
	I105x = 6320;
	I106x = 7950;
	I107x = -2846;
	I108x = 3383;
	I109x = -3418;
	I110x = -1556;
	I111x = 3474;
	I112x = -3208;
	I113x = 1451;
	I114x = -7134;
	I115x = -6424;
	I116x = -2016;
	I117x = 6185;
	I118x = 7761;
	I119x = 422;
	I120x = -2321;
	I121x = -3074;
	I122x = -7290;
	I123x = -3647;
	I124x = -2313;
	I125x = -7386;
	I126x = -2547;
	I127x = 2166;
	I128x = -1974;
	I129x = -946;
	I130x = -2723;
	I131x = 8187;
	I132x = -2435;
	I133x = -3721;
	I134x = -7294;
	I135x = -2908;
	I136x = -7564;
	I137x = 7103;
	I138x = 3192;
	I139x = 6020;
	I140x = -4797;
	I141x = 6724;
	I142x = -1737;
	I143x = -7281;
	I144x = 2350;
	I145x = 5886;
	I146x = 902;
	I147x = 6671;
	I148x = -2820;
	I149x = 4021;
	I150x = -4012;
	I151x = -775;
	I152x = -4677;
	I153x = 3219;
	I154x = -6646;
	I155x = 3772;
	I156x = -6106;
	I157x = -6077;
	I158x = 1361;
	I159x = 6774;
	I160x = 4298;
	I161x = 228;
	I162x = -3392;
	I163x = 1034;
	I164x = -1393;
	I165x = -3766;
	I166x = -5686;
	I167x = -3672;
	I168x = -6040;
	I169x = 6267;
	I170x = 2813;
	I171x = 5260;
	I172x = 7210;
	I173x = -4167;
	I174x = 2904;
	I175x = -1836;
	I176x = 7736;
	I177x = 5923;
	I178x = -1300;
	I179x = 3992;
	I180x = 6545;
	I181x = 2947;
	I182x = -3580;
	I183x = 7809;
	I184x = 2524;
	I185x = 494;
	I186x = 656;
	end
endmodule
[1.57347767 0.         0.         0.8235252  0.        ] 

 [12889, 0, 0, 6746, 0] 

 ['0011001001011001', '0000000000000000', '0000000000000000', '0001101001011010', '0000000000000000']
