module rom_input(EN,I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x);
	input EN;
	output [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
	reg [15:0]I0x,I1x,I2x,I3x,I4x,I5x,I6x,I7x,I8x,I9x,I10x,I11x,I12x,I13x,I14x,I15x,I16x,I17x,I18x,I19x,I20x,I21x,I22x,I23x,I24x,I25x,I26x,I27x,I28x,I29x,I30x,I31x,I32x,I33x,I34x,I35x,I36x,I37x,I38x,I39x,I40x,I41x,I42x,I43x,I44x,I45x,I46x,I47x,I48x,I49x,I50x,I51x,I52x,I53x,I54x,I55x,I56x,I57x,I58x,I59x,I60x,I61x,I62x,I63x,I64x,I65x,I66x,I67x,I68x,I69x,I70x,I71x,I72x,I73x,I74x,I75x,I76x,I77x,I78x,I79x,I80x,I81x,I82x,I83x,I84x,I85x,I86x,I87x,I88x,I89x,I90x,I91x,I92x,I93x,I94x,I95x,I96x,I97x,I98x,I99x,I100x,I101x,I102x,I103x,I104x,I105x,I106x,I107x,I108x,I109x,I110x,I111x,I112x,I113x,I114x,I115x,I116x,I117x,I118x,I119x,I120x,I121x,I122x,I123x,I124x,I125x,I126x,I127x,I128x,I129x,I130x,I131x,I132x,I133x,I134x,I135x,I136x,I137x,I138x,I139x,I140x,I141x,I142x,I143x,I144x,I145x,I146x,I147x,I148x,I149x,I150x,I151x,I152x,I153x,I154x,I155x,I156x,I157x,I158x,I159x,I160x,I161x,I162x,I163x,I164x,I165x,I166x,I167x,I168x,I169x,I170x,I171x,I172x,I173x,I174x,I175x,I176x,I177x,I178x,I179x,I180x,I181x,I182x,I183x,I184x,I185x,I186x;
always@(EN)
	begin
	I0x = 13;
	I1x = -12;
	I2x = -20;
	I3x = 18;
	I4x = 0;
	I5x = 7;
	I6x = -20;
	I7x = 8;
	I8x = -16;
	I9x = -23;
	I10x = -1;
	I11x = -28;
	I12x = 19;
	I13x = -5;
	I14x = 26;
	I15x = -26;
	I16x = 16;
	I17x = -22;
	I18x = 28;
	I19x = 23;
	I20x = 28;
	I21x = 22;
	I22x = 1;
	I23x = -29;
	I24x = -18;
	I25x = -20;
	I26x = -18;
	I27x = 31;
	I28x = -1;
	I29x = 28;
	I30x = 25;
	I31x = -7;
	I32x = 14;
	I33x = -25;
	I34x = 3;
	I35x = 23;
	I36x = 0;
	I37x = -30;
	I38x = 5;
	I39x = 14;
	I40x = -29;
	I41x = -9;
	I42x = -15;
	I43x = -21;
	I44x = 1;
	I45x = 28;
	I46x = 25;
	I47x = 25;
	I48x = -24;
	I49x = -20;
	I50x = 21;
	I51x = 0;
	I52x = -30;
	I53x = -24;
	I54x = -28;
	I55x = 11;
	I56x = -29;
	I57x = 6;
	I58x = -6;
	I59x = 29;
	I60x = 21;
	I61x = -23;
	I62x = -26;
	I63x = -13;
	I64x = -17;
	I65x = -11;
	I66x = 22;
	I67x = -1;
	I68x = 5;
	I69x = 0;
	I70x = -16;
	I71x = 22;
	I72x = 20;
	I73x = -17;
	I74x = 9;
	I75x = 8;
	I76x = -7;
	I77x = 14;
	I78x = -24;
	I79x = 21;
	I80x = -11;
	I81x = 0;
	I82x = 1;
	I83x = -26;
	I84x = -30;
	I85x = 8;
	I86x = -13;
	I87x = 5;
	I88x = 25;
	I89x = -27;
	I90x = 12;
	I91x = 27;
	I92x = -24;
	I93x = -3;
	I94x = 16;
	I95x = 0;
	I96x = 8;
	I97x = 2;
	I98x = 11;
	I99x = 0;
	I100x = 11;
	I101x = -24;
	I102x = 9;
	I103x = 18;
	I104x = 15;
	I105x = -28;
	I106x = -16;
	I107x = -19;
	I108x = -19;
	I109x = -5;
	I110x = -7;
	I111x = -25;
	I112x = -16;
	I113x = -22;
	I114x = -23;
	I115x = -4;
	I116x = 8;
	I117x = 25;
	I118x = 18;
	I119x = -19;
	I120x = 17;
	I121x = 15;
	I122x = -27;
	I123x = -24;
	I124x = 31;
	I125x = 2;
	I126x = -24;
	I127x = 10;
	I128x = -21;
	I129x = 0;
	I130x = -1;
	I131x = 20;
	I132x = 20;
	I133x = 22;
	I134x = -28;
	I135x = 25;
	I136x = 12;
	I137x = 19;
	I138x = -25;
	I139x = 4;
	I140x = -28;
	I141x = -14;
	I142x = 4;
	I143x = -5;
	I144x = -8;
	I145x = -17;
	I146x = 19;
	I147x = -21;
	I148x = -9;
	I149x = -20;
	I150x = -21;
	I151x = -3;
	I152x = -21;
	I153x = -19;
	I154x = 18;
	I155x = -21;
	I156x = -13;
	I157x = 19;
	I158x = 14;
	I159x = 1;
	I160x = -13;
	I161x = -4;
	I162x = 12;
	I163x = -16;
	I164x = 18;
	I165x = 0;
	I166x = -17;
	I167x = -29;
	I168x = -18;
	I169x = -25;
	I170x = 14;
	I171x = 27;
	I172x = -3;
	I173x = -31;
	I174x = 28;
	I175x = -8;
	I176x = -3;
	I177x = 14;
	I178x = 30;
	I179x = 9;
	I180x = 31;
	I181x = 8;
	I182x = -15;
	I183x = 2;
	I184x = 28;
	I185x = 10;
	I186x = -29;
	end
endmodule
[1.02887631 0.         2.46579106 1.25891637 1.42383812] 

 [32, 0, 78, 40, 45] 

 ['00100000', '00000000', '01001110', '00101000', '00101101']
